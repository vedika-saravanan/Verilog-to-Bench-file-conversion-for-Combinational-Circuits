module c7552 (N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, B241, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342);
input N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382;
output B241, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342;
wire N467, N469, N494, N528, N575, N578, N585, N590, N593, N596, N599, N604, N609, N614, N625, N628, N632, N636, N641, N642, N644, N651, N657, N660, N666, N672, N673, N674, N676, N682, N688, N689, N695, N700, N705, N706, N708, N715, N721, N727, N733, N734, N742, N748, N749, N750, N758, N759, N762, N768, N774, N780, N786, N794, N800, N806, N812, N814, N821, N827, N833, N839, N845, N853, N859, N865, N871, N886, N887, N957, N1028, N1029, N1109, N1115, N1116, N1119, N1125, N1132, N1136, N1141, N1147, N1154, N1160, N1167, N1174, N1175, N1182, N1189, N1194, N1199, N1206, N1211, N1218, N1222, N1227, N1233, N1240, N1244, N1249, N1256, N1263, N1270, N1277, N1284, N1287, N1290, N1293, N1296, N1299, N1302, N1305, N1308, N1311, N1314, N1317, N1320, N1323, N1326, N1329, N1332, N1335, N1338, N1341, N1344, N1347, N1350, N1353, N1356, N1359, N1362, N1365, N1368, N1371, N1374, N1377, N1380, N1383, N1386, N1389, N1392, N1395, N1398, N1401, N1404, N1407, N1410, N1413, N1416, N1419, N1422, N1425, N1428, N1431, N1434, N1437, N1440, N1443, N1446, N1449, N1452, N1455, N1458, N1461, N1464, N1467, N1470, N1473, N1476, N1479, N1482, N1485, N1537, N1551, N1649, N1703, N1708, N1713, N1721, N1758, N1782, N1783, N1789, N1793, N1794, N1795, N1796, N1797, N1798, N1799, N1805, N1811, N1812, N1813, N1814, N1815, N1816, N1817, N1818, N1819, N1820, N1821, N1822, N1828, N1829, N1830, N1832, N1833, N1834, N1835, N1839, N1840, N1841, N1842, N1843, N1845, N1851, N1857, N1858, N1859, N1860, N1861, N1862, N1863, N1864, N1865, N1866, N1867, N1868, N1869, N1870, N1871, N1872, N1873, N1874, N1875, N1876, N1877, N1878, N1879, N1880, N1881, N1882, N1883, N1884, N1885, N1892, N1899, N1906, N1913, N1919, N1926, N1927, N1928, N1929, N1930, N1931, N1932, N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942, N1943, N1944, N1945, N1946, N1947, N1953, N1957, N1958, N1959, N1960, N1961, N1962, N1963, N1965, N1966, N1967, N1968, N1969, N1970, N1971, N1972, N1973, N1974, N1975, N1976, N1977, N1983, N1989, N1990, N1991, N1992, N1993, N1994, N1995, N1996, N1997, N2003, N2010, N2011, N2012, N2013, N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024, N2031, N2038, N2045, N2052, N2058, N2064, N2065, N2066, N2067, N2068, N2069, N2070, N2071, N2072, N2073, N2074, N2081, N2086, N2107, N2108, N2110, N2111, N2112, N2113, N2114, N2115, N2117, N2171, N2172, N2230, N2231, N2235, N2239, N2240, N2241, N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249, N2250, N2251, N2252, N2253, N2254, N2255, N2256, N2257, N2267, N2268, N2269, N2274, N2275, N2277, N2278, N2279, N2280, N2281, N2282, N2283, N2284, N2285, N2286, N2287, N2293, N2299, N2300, N2301, N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2309, N2315, N2321, N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329, N2330, N2331, N2337, N2338, N2339, N2340, N2341, N2342, N2343, N2344, N2345, N2346, N2347, N2348, N2349, N2350, N2351, N2352, N2353, N2354, N2355, N2356, N2357, N2358, N2359, N2360, N2361, N2362, N2363, N2364, N2365, N2366, N2367, N2368, N2374, N2375, N2376, N2377, N2378, N2379, N2380, N2381, N2382, N2383, N2384, N2390, N2396, N2397, N2398, N2399, N2400, N2401, N2402, N2403, N2404, N2405, N2406, N2412, N2418, N2419, N2420, N2421, N2422, N2423, N2424, N2425, N2426, N2427, N2428, N2429, N2430, N2431, N2432, N2433, N2434, N2435, N2436, N2437, N2441, N2442, N2446, N2450, N2454, N2458, N2462, N2466, N2470, N2474, N2478, N2482, N2488, N2496, N2502, N2508, N2523, N2533, N2537, N2538, N2542, N2546, N2550, N2554, N2561, N2567, N2573, N2604, N2607, N2611, N2615, N2619, N2626, N2632, N2638, N2644, N2650, N2653, N2654, N2658, N2662, N2666, N2670, N2674, N2680, N2688, N2692, N2696, N2700, N2704, N2728, N2729, N2733, N2737, N2741, N2745, N2749, N2753, N2757, N2761, N2765, N2766, N2769, N2772, N2775, N2778, N2781, N2784, N2787, N2790, N2793, N2796, N2866, N2867, N2868, N2869, N2878, N2913, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N2988, N3005, N3006, N3007, N3008, N3009, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3032, N3033, N3034, N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3061, N3064, N3067, N3070, N3073, N3080, N3096, N3097, N3101, N3107, N3114, N3122, N3126, N3130, N3131, N3134, N3135, N3136, N3137, N3140, N3144, N3149, N3155, N3159, N3167, N3168, N3169, N3173, N3178, N3184, N3185, N3189, N3195, N3202, N3210, N3211, N3215, N3221, N3228, N3229, N3232, N3236, N3241, N3247, N3251, N3255, N3259, N3263, N3267, N3273, N3281, N3287, N3293, N3299, N3303, N3307, N3311, N3315, N3322, N3328, N3334, N3340, N3343, N3349, N3355, N3361, N3362, N3363, N3364, N3365, N3366, N3367, N3368, N3369, N3370, N3371, N3372, N3373, N3374, N3375, N3379, N3380, N3381, N3384, N3390, N3398, N3404, N3410, N3416, N3420, N3424, N3428, N3432, N3436, N3440, N3444, N3448, N3452, N3453, N3454, N3458, N3462, N3466, N3470, N3474, N3478, N3482, N3486, N3487, N3490, N3493, N3496, N3499, N3502, N3507, N3510, N3515, N3518, N3521, N3524, N3527, N3530, N3535, N3539, N3542, N3545, N3548, N3551, N3552, N3553, N3557, N3560, N3563, N3566, N3569, N3570, N3571, N3574, N3577, N3580, N3583, N3586, N3589, N3592, N3595, N3598, N3601, N3604, N3607, N3610, N3613, N3616, N3619, N3622, N3625, N3628, N3631, N3634, N3637, N3640, N3643, N3646, N3649, N3652, N3655, N3658, N3661, N3664, N3667, N3670, N3673, N3676, N3679, N3682, N3685, N3688, N3691, N3694, N3697, N3700, N3703, N3706, N3709, N3712, N3715, N3718, N3721, N3724, N3727, N3730, N3733, N3736, N3739, N3742, N3745, N3748, N3751, N3754, N3757, N3760, N3763, N3766, N3769, N3772, N3775, N3778, N3781, N3782, N3783, N3786, N3789, N3792, N3795, N3798, N3801, N3804, N3807, N3810, N3813, N3816, N3819, N3822, N3825, N3828, N3831, N3834, N3837, N3840, N3843, N3846, N3849, N3852, N3855, N3858, N3861, N3864, N3867, N3870, N3873, N3876, N3879, N3882, N3885, N3888, N3891, N3953, N3954, N3955, N3956, N3958, N3964, N4193, N4303, N4308, N4313, N4326, N4327, N4333, N4334, N4411, N4412, N4463, N4464, N4465, N4466, N4467, N4468, N4469, N4470, N4471, N4472, N4473, N4474, N4475, N4476, N4477, N4478, N4479, N4480, N4481, N4482, N4483, N4484, N4485, N4486, N4487, N4488, N4489, N4490, N4491, N4492, N4493, N4494, N4495, N4496, N4497, N4498, N4499, N4500, N4501, N4502, N4503, N4504, N4505, N4506, N4507, N4508, N4509, N4510, N4511, N4512, N4513, N4514, N4515, N4516, N4517, N4518, N4519, N4520, N4521, N4522, N4523, N4524, N4525, N4526, N4527, N4528, N4529, N4530, N4531, N4532, N4533, N4534, N4535, N4536, N4537, N4538, N4539, N4540, N4541, N4542, N4543, N4544, N4545, N4549, N4555, N4562, N4563, N4566, N4570, N4575, N4576, N4577, N4581, N4586, N4592, N4593, N4597, N4603, N4610, N4611, N4612, N4613, N4614, N4615, N4616, N4617, N4618, N4619, N4620, N4621, N4622, N4623, N4624, N4625, N4626, N4627, N4628, N4629, N4630, N4631, N4632, N4633, N4634, N4635, N4636, N4637, N4638, N4639, N4640, N4641, N4642, N4643, N4644, N4645, N4646, N4647, N4648, N4649, N4650, N4651, N4652, N4653, N4656, N4657, N4661, N4667, N4674, N4675, N4678, N4682, N4687, N4693, N4694, N4695, N4696, N4697, N4698, N4699, N4700, N4701, N4702, N4706, N4711, N4717, N4718, N4722, N4728, N4735, N4743, N4744, N4745, N4746, N4747, N4748, N4749, N4750, N4751, N4752, N4753, N4754, N4755, N4756, N4757, N4758, N4759, N4760, N4761, N4762, N4763, N4764, N4765, N4766, N4767, N4768, N4769, N4775, N4776, N4777, N4778, N4779, N4780, N4781, N4782, N4783, N4784, N4789, N4790, N4793, N4794, N4795, N4796, N4799, N4800, N4801, N4802, N4803, N4806, N4809, N4810, N4813, N4814, N4817, N4820, N4823, N4826, N4829, N4832, N4835, N4838, N4841, N4844, N4847, N4850, N4853, N4856, N4859, N4862, N4865, N4868, N4871, N4874, N4877, N4880, N4883, N4886, N4889, N4892, N4895, N4898, N4901, N4904, N4907, N4910, N4913, N4916, N4919, N4922, N4925, N4928, N4931, N4934, N4937, N4940, N4943, N4946, N4949, N4952, N4955, N4958, N4961, N4964, N4967, N4970, N4973, N4976, N4979, N4982, N4985, N4988, N4991, N4994, N4997, N5000, N5003, N5006, N5009, N5012, N5015, N5018, N5021, N5024, N5027, N5030, N5033, N5036, N5039, N5042, N5045, N5046, N5047, N5048, N5049, N5052, N5055, N5058, N5061, N5064, N5065, N5066, N5067, N5068, N5071, N5074, N5077, N5080, N5083, N5086, N5089, N5092, N5095, N5098, N5101, N5104, N5107, N5110, N5111, N5112, N5113, N5114, N5117, N5120, N5123, N5126, N5129, N5132, N5135, N5138, N5141, N5144, N5147, N5150, N5153, N5156, N5159, N5162, N5165, N5166, N5167, N5168, N5169, N5170, N5171, N5172, N5173, N5174, N5175, N5176, N5177, N5178, N5179, N5180, N5181, N5182, N5183, N5184, N5185, N5186, N5187, N5188, N5189, N5190, N5191, N5192, N5193, N5196, N5197, N5198, N5199, N5200, N5201, N5202, N5203, N5204, N5205, N5206, N5207, N5208, N5209, N5210, N5211, N5212, N5213, N5283, N5284, N5285, N5286, N5287, N5288, N5289, N5290, N5291, N5292, N5293, N5294, N5295, N5296, N5297, N5298, N5299, N5300, N5314, N5315, N5316, N5317, N5318, N5319, N5320, N5321, N5322, N5323, N5324, N5363, N5364, N5365, N5366, N5367, N5425, N5426, N5427, N5429, N5430, N5431, N5432, N5433, N5451, N5452, N5453, N5454, N5455, N5456, N5457, N5469, N5474, N5475, N5476, N5477, N5571, N5572, N5573, N5574, N5584, N5585, N5586, N5587, N5602, N5603, N5604, N5605, N5631, N5632, N5640, N5654, N5670, N5683, N5690, N5697, N5707, N5718, N5728, N5735, N5736, N5740, N5744, N5747, N5751, N5755, N5758, N5762, N5766, N5769, N5770, N5771, N5778, N5789, N5799, N5807, N5821, N5837, N5850, N5856, N5863, N5870, N5881, N5892, N5898, N5905, N5915, N5926, N5936, N5943, N5944, N5945, N5946, N5947, N5948, N5949, N5950, N5951, N5952, N5953, N5954, N5955, N5956, N5957, N5958, N5959, N5960, N5966, N5967, N5968, N5969, N5970, N5971, N5972, N5973, N5974, N5975, N5976, N5977, N5978, N5979, N5980, N5981, N5989, N5990, N5991, N5996, N6000, N6003, N6009, N6014, N6018, N6021, N6022, N6023, N6024, N6025, N6026, N6027, N6028, N6029, N6030, N6031, N6032, N6033, N6034, N6035, N6036, N6037, N6038, N6039, N6040, N6041, N6047, N6052, N6056, N6059, N6060, N6061, N6062, N6063, N6064, N6065, N6066, N6067, N6068, N6069, N6070, N6071, N6072, N6073, N6074, N6075, N6076, N6077, N6078, N6079, N6083, N6087, N6090, N6091, N6092, N6093, N6094, N6095, N6096, N6097, N6098, N6099, N6100, N6101, N6102, N6103, N6104, N6105, N6106, N6107, N6108, N6109, N6110, N6111, N6112, N6113, N6114, N6115, N6116, N6117, N6118, N6119, N6120, N6121, N6122, N6123, N6124, N6125, N6126, N6127, N6131, N6135, N6136, N6137, N6141, N6145, N6148, N6149, N6150, N6151, N6152, N6153, N6154, N6155, N6156, N6157, N6158, N6159, N6160, N6161, N6162, N6163, N6164, N6165, N6166, N6170, N6174, N6177, N6181, N6182, N6183, N6184, N6185, N6186, N6187, N6188, N6189, N6190, N6191, N6192, N6193, N6194, N6195, N6196, N6199, N6202, N6203, N6204, N6207, N6210, N6213, N6214, N6217, N6220, N6223, N6224, N6225, N6226, N6227, N6228, N6229, N6230, N6231, N6232, N6235, N6236, N6239, N6240, N6241, N6242, N6243, N6246, N6249, N6252, N6255, N6256, N6257, N6258, N6259, N6260, N6261, N6262, N6263, N6266, N6540, N6541, N6542, N6543, N6544, N6545, N6546, N6547, N6555, N6556, N6557, N6558, N6559, N6560, N6561, N6569, N6594, N6595, N6596, N6597, N6598, N6599, N6600, N6601, N6602, N6603, N6604, N6605, N6606, N6621, N6622, N6623, N6624, N6625, N6626, N6627, N6628, N6629, N6639, N6640, N6641, N6642, N6643, N6644, N6645, N6646, N6647, N6648, N6649, N6650, N6651, N6652, N6653, N6654, N6655, N6656, N6657, N6658, N6659, N6660, N6661, N6668, N6677, N6678, N6679, N6680, N6681, N6682, N6683, N6684, N6685, N6686, N6687, N6688, N6689, N6690, N6702, N6703, N6704, N6705, N6706, N6707, N6708, N6709, N6710, N6711, N6712, N6729, N6730, N6731, N6732, N6733, N6734, N6735, N6736, N6741, N6742, N6743, N6744, N6751, N6752, N6753, N6754, N6755, N6756, N6757, N6758, N6761, N6762, N6766, N6767, N6768, N6769, N6770, N6771, N6772, N6773, N6774, N6775, N6776, N6777, N6778, N6779, N6780, N6781, N6782, N6783, N6784, N6787, N6788, N6789, N6790, N6791, N6792, N6793, N6794, N6795, N6796, N6797, N6800, N6803, N6806, N6809, N6812, N6815, N6818, N6821, N6824, N6827, N6830, N6833, N6836, N6837, N6838, N6839, N6840, N6841, N6842, N6843, N6844, N6845, N6848, N6849, N6850, N6851, N6852, N6853, N6854, N6855, N6856, N6857, N6858, N6859, N6860, N6861, N6862, N6863, N6864, N6865, N6866, N6867, N6870, N6871, N6872, N6873, N6874, N6875, N6876, N6877, N6878, N6879, N6880, N6881, N6884, N6885, N6886, N6887, N6888, N6889, N6890, N6891, N6892, N6893, N6894, N6901, N6912, N6923, N6929, N6936, N6946, N6957, N6967, N6968, N6969, N6970, N6977, N6988, N6998, N7006, N7020, N7036, N7049, N7055, N7056, N7057, N7060, N7061, N7062, N7063, N7064, N7065, N7066, N7067, N7068, N7073, N7077, N7080, N7086, N7091, N7095, N7098, N7099, N7100, N7103, N7104, N7105, N7106, N7107, N7114, N7125, N7136, N7142, N7149, N7159, N7170, N7180, N7187, N7188, N7191, N7194, N7198, N7202, N7205, N7209, N7213, N7216, N7219, N7222, N7229, N7240, N7250, N7258, N7272, N7288, N7301, N7307, N7314, N7318, N7322, N7325, N7328, N7331, N7334, N7337, N7340, N7343, N7346, N7351, N7355, N7358, N7364, N7369, N7373, N7376, N7377, N7378, N7381, N7384, N7387, N7391, N7394, N7398, N7402, N7405, N7408, N7411, N7414, N7417, N7420, N7423, N7426, N7429, N7432, N7435, N7438, N7441, N7444, N7447, N7450, N7453, N7456, N7459, N7462, N7465, N7468, N7471, N7474, N7477, N7478, N7479, N7482, N7485, N7488, N7491, N7494, N7497, N7500, N7503, N7506, N7509, N7512, N7515, N7518, N7521, N7524, N7527, N7530, N7533, N7536, N7539, N7542, N7545, N7548, N7551, N7552, N7553, N7556, N7557, N7558, N7559, N7560, N7563, N7566, N7569, N7572, N7573, N7574, N7577, N7580, N7581, N7582, N7585, N7588, N7591, N7609, N7613, N7620, N7649, N7650, N7655, N7659, N7668, N7671, N7744, N7822, N7825, N7826, N7852, N8114, N8117, N8131, N8134, N8144, N8145, N8146, N8156, N8166, N8169, N8183, N8186, N8196, N8200, N8204, N8208, N8216, N8217, N8218, N8219, N8232, N8233, N8242, N8243, N8244, N8245, N8246, N8247, N8248, N8249, N8250, N8251, N8252, N8253, N8254, N8260, N8261, N8262, N8269, N8274, N8275, N8276, N8277, N8278, N8279, N8280, N8281, N8282, N8283, N8284, N8285, N8288, N8294, N8295, N8296, N8297, N8298, N8307, N8315, N8317, N8319, N8321, N8322, N8323, N8324, N8325, N8326, N8333, N8337, N8338, N8339, N8340, N8341, N8342, N8343, N8344, N8345, N8346, N8347, N8348, N8349, N8350, N8351, N8352, N8353, N8354, N8355, N8356, N8357, N8358, N8365, N8369, N8370, N8371, N8372, N8373, N8374, N8375, N8376, N8377, N8378, N8379, N8380, N8381, N8382, N8383, N8384, N8385, N8386, N8387, N8388, N8389, N8390, N8391, N8392, N8393, N8394, N8404, N8405, N8409, N8410, N8411, N8412, N8415, N8416, N8417, N8418, N8421, N8430, N8433, N8434, N8435, N8436, N8437, N8438, N8439, N8440, N8441, N8442, N8443, N8444, N8447, N8448, N8449, N8450, N8451, N8452, N8453, N8454, N8455, N8456, N8457, N8460, N8463, N8466, N8469, N8470, N8471, N8474, N8477, N8480, N8483, N8484, N8485, N8488, N8489, N8490, N8491, N8492, N8493, N8494, N8495, N8496, N8497, N8500, N8501, N8502, N8503, N8504, N8505, N8506, N8507, N8508, N8509, N8510, N8511, N8512, N8513, N8514, N8515, N8516, N8517, N8518, N8519, N8522, N8525, N8528, N8531, N8534, N8537, N8538, N8539, N8540, N8541, N8545, N8546, N8547, N8548, N8551, N8552, N8553, N8554, N8555, N8558, N8561, N8564, N8565, N8566, N8569, N8572, N8575, N8578, N8579, N8580, N8583, N8586, N8589, N8592, N8595, N8598, N8601, N8604, N8607, N8608, N8609, N8610, N8615, N8616, N8617, N8618, N8619, N8624, N8625, N8626, N8627, N8632, N8633, N8634, N8637, N8638, N8639, N8644, N8645, N8646, N8647, N8648, N8653, N8654, N8655, N8660, N8663, N8666, N8669, N8672, N8675, N8678, N8681, N8684, N8687, N8690, N8693, N8696, N8699, N8702, N8705, N8708, N8711, N8714, N8717, N8718, N8721, N8724, N8727, N8730, N8733, N8734, N8735, N8738, N8741, N8744, N8747, N8750, N8753, N8754, N8755, N8756, N8757, N8760, N8763, N8766, N8769, N8772, N8775, N8778, N8781, N8784, N8787, N8790, N8793, N8796, N8799, N8802, N8805, N8808, N8811, N8814, N8815, N8816, N8817, N8818, N8840, N8857, N8861, N8862, N8863, N8864, N8865, N8866, N8871, N8874, N8878, N8879, N8880, N8881, N8882, N8883, N8884, N8885, N8886, N8887, N8888, N8898, N8902, N8920, N8924, N8927, N8931, N8943, N8950, N8956, N8959, N8960, N8963, N8966, N8991, N8992, N8995, N8996, N9001, N9005, N9024, N9025, N9029, N9035, N9053, N9054, N9064, N9065, N9066, N9067, N9068, N9071, N9072, N9073, N9074, N9077, N9079, N9082, N9083, N9086, N9087, N9088, N9089, N9092, N9093, N9094, N9095, N9098, N9099, N9103, N9107, N9111, N9117, N9127, N9146, N9149, N9159, N9160, N9161, N9165, N9169, N9173, N9179, N9180, N9181, N9182, N9183, N9193, N9203, N9206, N9220, N9223, N9234, N9235, N9236, N9237, N9238, N9242, N9243, N9244, N9245, N9246, N9247, N9248, N9249, N9250, N9251, N9252, N9256, N9257, N9258, N9259, N9260, N9261, N9262, N9265, N9268, N9271, N9272, N9273, N9274, N9275, N9276, N9280, N9285, N9286, N9287, N9288, N9290, N9292, N9294, N9296, N9297, N9298, N9299, N9300, N9301, N9307, N9314, N9315, N9318, N9319, N9320, N9321, N9322, N9323, N9324, N9326, N9332, N9339, N9344, N9352, N9354, N9356, N9358, N9359, N9360, N9361, N9362, N9363, N9364, N9365, N9366, N9367, N9368, N9369, N9370, N9371, N9372, N9375, N9381, N9382, N9383, N9384, N9385, N9392, N9393, N9394, N9395, N9396, N9397, N9398, N9399, N9400, N9401, N9402, N9407, N9408, N9412, N9413, N9414, N9415, N9416, N9417, N9418, N9419, N9420, N9421, N9422, N9423, N9426, N9429, N9432, N9435, N9442, N9445, N9454, N9455, N9456, N9459, N9460, N9461, N9462, N9465, N9466, N9467, N9468, N9473, N9476, N9477, N9478, N9485, N9488, N9493, N9494, N9495, N9498, N9499, N9500, N9505, N9506, N9507, N9508, N9509, N9514, N9515, N9516, N9517, N9520, N9526, N9531, N9539, N9540, N9541, N9543, N9551, N9555, N9556, N9557, N9560, N9561, N9562, N9563, N9564, N9565, N9566, N9567, N9568, N9569, N9570, N9571, N9575, N9579, N9581, N9582, N9585, N9591, N9592, N9593, N9594, N9595, N9596, N9597, N9598, N9599, N9600, N9601, N9602, N9603, N9604, N9605, N9608, N9611, N9612, N9613, N9614, N9615, N9616, N9617, N9618, N9621, N9622, N9623, N9624, N9626, N9629, N9632, N9635, N9642, N9645, N9646, N9649, N9650, N9653, N9656, N9659, N9660, N9661, N9662, N9663, N9666, N9667, N9670, N9671, N9674, N9675, N9678, N9679, N9682, N9685, N9690, N9691, N9692, N9695, N9698, N9702, N9707, N9710, N9711, N9714, N9715, N9716, N9717, N9720, N9721, N9722, N9723, N9726, N9727, N9732, N9733, N9734, N9735, N9736, N9737, N9738, N9739, N9740, N9741, N9742, N9754, N9758, N9762, N9763, N9764, N9765, N9766, N9767, N9768, N9769, N9773, N9774, N9775, N9779, N9784, N9785, N9786, N9790, N9791, N9795, N9796, N9797, N9798, N9799, N9800, N9801, N9802, N9803, N9805, N9806, N9809, N9813, N9814, N9815, N9816, N9817, N9820, N9825, N9826, N9827, N9828, N9829, N9830, N9835, N9836, N9837, N9838, N9846, N9847, N9862, N9863, N9866, N9873, N9876, N9890, N9891, N9892, N9893, N9894, N9895, N9896, N9897, N9898, N9899, N9900, N9901, N9902, N9903, N9904, N9905, N9906, N9907, N9908, N9909, N9910, N9911, N9917, N9923, N9924, N9925, N9932, N9935, N9938, N9939, N9945, N9946, N9947, N9948, N9949, N9953, N9954, N9955, N9956, N9957, N9958, N9959, N9960, N9961, N9964, N9967, N9968, N9969, N9970, N9971, N9972, N9973, N9974, N9975, N9976, N9977, N9978, N9979, N9982, N9983, N9986, N9989, N9992, N9995, N9996, N9997, N9998, N9999, N10002, N10003, N10006, N10007, N10010, N10013, N10014, N10015, N10016, N10017, N10018, N10019, N10020, N10021, N10022, N10023, N10024, N10026, N10028, N10032, N10033, N10034, N10035, N10036, N10037, N10038, N10039, N10040, N10041, N10042, N10043, N10050, N10053, N10054, N10055, N10056, N10057, N10058, N10059, N10060, N10061, N10062, N10067, N10070, N10073, N10076, N10077, N10082, N10083, N10084, N10085, N10086, N10093, N10094, N10105, N10106, N10107, N10108, N10113, N10114, N10115, N10116, N10119, N10124, N10130, N10131, N10132, N10133, N10134, N10135, N10136, N10137, N10138, N10139, N10140, N10141, N10148, N10155, N10156, N10157, N10158, N10159, N10160, N10161, N10162, N10163, N10164, N10165, N10170, N10173, N10176, N10177, N10178, N10179, N10180, N10183, N10186, N10189, N10192, N10195, N10196, N10197, N10200, N10203, N10204, N10205, N10206, N10212, N10213, N10230, N10231, N10232, N10233, N10234, N10237, N10238, N10239, N10240, N10241, N10242, N10247, N10248, N10259, N10264, N10265, N10266, N10267, N10268, N10269, N10270, N10271, N10272, N10273, N10278, N10279, N10280, N10281, N10282, N10283, N10287, N10288, N10289, N10290, N10291, N10292, N10293, N10294, N10295, N10296, N10299, N10300, N10301, N10306, N10307, N10308, N10311, N10314, N10315, N10316, N10317, N10318, N10321, N10324, N10325, N10326, N10327, N10328, N10329, N10330, N10331, N10332, N10333, N10334, N10337, N10338, N10339, N10340, N10341, N10344, N10354, N10357, N10360, N10367, N10375, N10381, N10388, N10391, N10399, N10402, N10406, N10409, N10412, N10415, N10419, N10422, N10425, N10428, N10431, N10432, N10437, N10438, N10439, N10440, N10441, N10444, N10445, N10450, N10451, N10455, N10456, N10465, N10466, N10479, N10497, N10509, N10512, N10515, N10516, N10517, N10518, N10519, N10522, N10525, N10528, N10531, N10534, N10535, N10536, N10539, N10542, N10543, N10544, N10545, N10546, N10547, N10548, N10549, N10550, N10551, N10552, N10553, N10554, N10555, N10556, N10557, N10558, N10559, N10560, N10561, N10562, N10563, N10564, N10565, N10566, N10567, N10568, N10569, N10570, N10571, N10572, N10573, N10577, N10581, N10582, N10583, N10587, N10588, N10589, N10594, N10595, N10596, N10597, N10598, N10602, N10609, N10610, N10621, N10626, N10627, N10629, N10631, N10637, N10638, N10639, N10640, N10642, N10643, N10644, N10645, N10647, N10648, N10649, N10652, N10659, N10662, N10665, N10668, N10671, N10672, N10673, N10674, N10675, N10678, N10681, N10682, N10683, N10684, N10685, N10686, N10687, N10688, N10689, N10690, N10691, N10694, N10695, N10696, N10697, N10698, N10701, N10705, N10707, N10708, N10709, N10710, N10719, N10720, N10730, N10731, N10737, N10738, N10739, N10746, N10747, N10748, N10749, N10750, N10753, N10754, N10764, N10765, N10766, N10767, N10768, N10769, N10770, N10771, N10772, N10773, N10774, N10775, N10776, N10778, N10781, N10784, N10789, N10792, N10796, N10797, N10798, N10799, N10800, N10803, N10806, N10809, N10812, N10815, N10816, N10817, N10820, N10823, N10824, N10825, N10826, N10832, N10833, N10834, N10835, N10836, N10845, N10846, N10857, N10862, N10863, N10864, N10865, N10866, N10867, N10872, N10873, N10874, N10875, N10876, N10879, N10882, N10883, N10884, N10885, N10886, N10887, N10888, N10889, N10890, N10891, N10892, N10895, N10896, N10897, N10898, N10899, N10902, N10909, N10910, N10915, N10916, N10917, N10918, N10919, N10922, N10923, N10928, N10931, N10934, N10935, N10936, N10937, N10938, N10941, N10944, N10947, N10950, N10953, N10954, N10955, N10958, N10961, N10962, N10963, N10964, N10969, N10970, N10981, N10986, N10987, N10988, N10989, N10990, N10991, N10992, N10995, N10998, N10999, N11000, N11001, N11002, N11003, N11004, N11005, N11006, N11007, N11008, N11011, N11012, N11013, N11014, N11015, N11018, N11023, N11024, N11027, N11028, N11029, N11030, N11031, N11034, N11035, N11040, N11041, N11042, N11043, N11044, N11047, N11050, N11053, N11056, N11059, N11062, N11065, N11066, N11067, N11070, N11073, N11074, N11075, N11076, N11077, N11078, N11095, N11098, N11099, N11100, N11103, N11106, N11107, N11108, N11109, N11110, N11111, N11112, N11113, N11114, N11115, N11116, N11117, N11118, N11119, N11120, N11121, N11122, N11123, N11124, N11127, N11130, N11137, N11138, N11139, N11140, N11141, N11142, N11143, N11144, N11145, N11152, N11153, N11154, N11155, N11156, N11159, N11162, N11165, N11168, N11171, N11174, N11177, N11180, N11183, N11184, N11185, N11186, N11187, N11188, N11205, N11210, N11211, N11212, N11213, N11214, N11215, N11216, N11217, N11218, N11219, N11220, N11222, N11223, N11224, N11225, N11226, N11227, N11228, N11229, N11231, N11232, N11233, N11236, N11239, N11242, N11243, N11244, N11245, N11246, N11250, N11252, N11257, N11260, N11261, N11262, N11263, N11264, N11265, N11267, N11268, N11269, N11270, N11272, N11277, N11278, N11279, N11280, N11282, N11283, N11284, N11285, N11286, N11288, N11289, N11290, N11291, N11292, N11293, N11294, N11295, N11296, N11297, N11298, N11299, N11302, N11307, N11308, N11309, N11312, N11313, N11314, N11315, N11316, N11317, N11320, N11321, N11323, N11327, N11328, N11329, N11331, N11335, N11336, N11337, N11338, N11339, N11341;

buff U1 (N387,N1);
buff U2 (N388,N1);
not U3 (N467,N57);
and U4 (N469,N134,N133);
buff U5 (N478,N248);
buff U6 (N482,N254);
buff U7 (N484,N257);
buff U8 (N486,N260);
buff U9 (N489,N263);
buff U10 (N492,N267);
and U11 (N494,N162,N172,N188,N199);
buff U12 (N501,N274);
buff U13 (N505,N280);
buff U14 (N507,N283);
buff U15 (N509,N286);
buff U16 (N511,N289);
buff U17 (N513,N293);
buff U18 (N515,N296);
buff U19 (N517,N299);
buff U20 (N519,N303);
and U21 (N528,N150,N184,N228,N240);
buff U22 (N535,N307);
buff U23 (N537,N310);
buff U24 (N539,N313);
buff U25 (N541,N316);
buff U26 (N543,N319);
buff U27 (N545,N322);
buff U28 (N547,N325);
buff U29 (N549,N328);
buff U30 (N551,N331);
buff U31 (N553,N334);
buff U32 (N556,N337);
buff U33 (N559,N343);
buff U34 (N561,N346);
buff U35 (N563,N349);
buff U36 (N565,N352);
buff U37 (N567,N355);
buff U38 (N569,N358);
buff U39 (N571,N361);
buff U40 (N573,N364);
and U41 (N575,N183,N182,N185,N186);
and U42 (N578,N210,N152,N218,N230);
not U43 (N582,N15);
not U44 (N585,N5);
buff U45 (N590,N1);
not U46 (N593,N5);
not U47 (N596,N5);
not U48 (N599,N289);
not U49 (N604,N299);
not U50 (N609,N303);
buff U51 (N614,N38);
buff U52 (N625,N15);
nand U53 (N628,N12,N9);
nand U54 (N632,N12,N9);
buff U55 (N636,N38);
not U56 (N641,N245);
not U57 (N642,N248);
buff U58 (N643,N251);
not U59 (N644,N251);
not U60 (N651,N254);
buff U61 (N657,N106);
not U62 (N660,N257);
not U63 (N666,N260);
not U64 (N672,N263);
not U65 (N673,N267);
not U66 (N674,N106);
buff U67 (N676,N18);
buff U68 (N682,N18);
and U69 (N688,N382,N263);
buff U70 (N689,N18);
not U71 (N695,N18);
nand U72 (N700,N382,N267);
not U73 (N705,N271);
not U74 (N706,N274);
buff U75 (N707,N277);
not U76 (N708,N277);
not U77 (N715,N280);
not U78 (N721,N283);
not U79 (N727,N286);
not U80 (N733,N289);
not U81 (N734,N293);
not U82 (N742,N296);
not U83 (N748,N299);
not U84 (N749,N303);
buff U85 (N750,N367);
not U86 (N758,N307);
not U87 (N759,N310);
not U88 (N762,N313);
not U89 (N768,N316);
not U90 (N774,N319);
not U91 (N780,N322);
not U92 (N786,N325);
not U93 (N794,N328);
not U94 (N800,N331);
not U95 (N806,N334);
not U96 (N812,N337);
buff U97 (N813,N340);
not U98 (N814,N340);
not U99 (N821,N343);
not U100 (N827,N346);
not U101 (N833,N349);
not U102 (N839,N352);
not U103 (N845,N355);
not U104 (N853,N358);
not U105 (N859,N361);
not U106 (N865,N364);
buff U107 (N871,N367);
nand U108 (N881,N467,N585);
not U109 (N882,N528);
not U110 (N883,N578);
not U111 (N884,N575);
not U112 (N885,N494);
and U113 (N886,N528,N578);
and U114 (N887,N575,N494);
buff U115 (N889,N590);
buff U116 (N945,N657);
not U117 (N957,N688);
and U118 (N1028,N382,N641);
nand U119 (N1029,N382,N705);
and U120 (N1109,N469,N596);
nand U121 (N1110,N242,N593);
not U122 (N1111,N625);
nand U123 (N1112,N242,N593);
nand U124 (N1113,N469,N596);
not U125 (N1114,N625);
not U126 (N1115,N871);
buff U127 (N1116,N590);
buff U128 (N1119,N628);
buff U129 (N1125,N682);
buff U130 (N1132,N628);
buff U131 (N1136,N682);
buff U132 (N1141,N628);
buff U133 (N1147,N682);
buff U134 (N1154,N632);
buff U135 (N1160,N676);
and U136 (N1167,N700,N614);
and U137 (N1174,N700,N614);
buff U138 (N1175,N682);
buff U139 (N1182,N676);
not U140 (N1189,N657);
not U141 (N1194,N676);
not U142 (N1199,N682);
not U143 (N1206,N689);
buff U144 (N1211,N695);
not U145 (N1218,N750);
not U146 (N1222,N1028);
buff U147 (N1227,N632);
buff U148 (N1233,N676);
buff U149 (N1240,N632);
buff U150 (N1244,N676);
buff U151 (N1249,N689);
buff U152 (N1256,N689);
buff U153 (N1263,N695);
buff U154 (N1270,N689);
buff U155 (N1277,N689);
buff U156 (N1284,N700);
buff U157 (N1287,N614);
buff U158 (N1290,N666);
buff U159 (N1293,N660);
buff U160 (N1296,N651);
buff U161 (N1299,N614);
buff U162 (N1302,N644);
buff U163 (N1305,N700);
buff U164 (N1308,N614);
buff U165 (N1311,N614);
buff U166 (N1314,N666);
buff U167 (N1317,N660);
buff U168 (N1320,N651);
buff U169 (N1323,N644);
buff U170 (N1326,N609);
buff U171 (N1329,N604);
buff U172 (N1332,N742);
buff U173 (N1335,N599);
buff U174 (N1338,N727);
buff U175 (N1341,N721);
buff U176 (N1344,N715);
buff U177 (N1347,N734);
buff U178 (N1350,N708);
buff U179 (N1353,N609);
buff U180 (N1356,N604);
buff U181 (N1359,N742);
buff U182 (N1362,N734);
buff U183 (N1365,N599);
buff U184 (N1368,N727);
buff U185 (N1371,N721);
buff U186 (N1374,N715);
buff U187 (N1377,N708);
buff U188 (N1380,N806);
buff U189 (N1383,N800);
buff U190 (N1386,N794);
buff U191 (N1389,N786);
buff U192 (N1392,N780);
buff U193 (N1395,N774);
buff U194 (N1398,N768);
buff U195 (N1401,N762);
buff U196 (N1404,N806);
buff U197 (N1407,N800);
buff U198 (N1410,N794);
buff U199 (N1413,N780);
buff U200 (N1416,N774);
buff U201 (N1419,N768);
buff U202 (N1422,N762);
buff U203 (N1425,N786);
buff U204 (N1428,N636);
buff U205 (N1431,N636);
buff U206 (N1434,N865);
buff U207 (N1437,N859);
buff U208 (N1440,N853);
buff U209 (N1443,N845);
buff U210 (N1446,N839);
buff U211 (N1449,N833);
buff U212 (N1452,N827);
buff U213 (N1455,N821);
buff U214 (N1458,N814);
buff U215 (N1461,N865);
buff U216 (N1464,N859);
buff U217 (N1467,N853);
buff U218 (N1470,N839);
buff U219 (N1473,N833);
buff U220 (N1476,N827);
buff U221 (N1479,N821);
buff U222 (N1482,N845);
buff U223 (N1485,N814);
not U224 (N1489,N1109);
buff U225 (N1490,N1116);
and U226 (N1537,N957,N614);
and U227 (N1551,N614,N957);
and U228 (N1649,N1029,N636);
buff U229 (N1703,N957);
nor U230 (N1708,N957,N614);
buff U231 (N1713,N957);
nor U232 (N1721,N614,N957);
buff U233 (N1758,N1029);
and U234 (N1781,N163,N1116);
and U235 (N1782,N170,N1125);
not U236 (N1783,N1125);
not U237 (N1789,N1136);
and U238 (N1793,N169,N1125);
and U239 (N1794,N168,N1125);
and U240 (N1795,N167,N1125);
and U241 (N1796,N166,N1136);
and U242 (N1797,N165,N1136);
and U243 (N1798,N164,N1136);
not U244 (N1799,N1147);
not U245 (N1805,N1160);
and U246 (N1811,N177,N1147);
and U247 (N1812,N176,N1147);
and U248 (N1813,N175,N1147);
and U249 (N1814,N174,N1147);
and U250 (N1815,N173,N1147);
and U251 (N1816,N157,N1160);
and U252 (N1817,N156,N1160);
and U253 (N1818,N155,N1160);
and U254 (N1819,N154,N1160);
and U255 (N1820,N153,N1160);
not U256 (N1821,N1284);
not U257 (N1822,N1287);
not U258 (N1828,N1290);
not U259 (N1829,N1293);
not U260 (N1830,N1296);
not U261 (N1832,N1299);
not U262 (N1833,N1302);
not U263 (N1834,N1305);
not U264 (N1835,N1308);
not U265 (N1839,N1311);
not U266 (N1840,N1314);
not U267 (N1841,N1317);
not U268 (N1842,N1320);
not U269 (N1843,N1323);
not U270 (N1845,N1175);
not U271 (N1851,N1182);
and U272 (N1857,N181,N1175);
and U273 (N1858,N171,N1175);
and U274 (N1859,N180,N1175);
and U275 (N1860,N179,N1175);
and U276 (N1861,N178,N1175);
and U277 (N1862,N161,N1182);
and U278 (N1863,N151,N1182);
and U279 (N1864,N160,N1182);
and U280 (N1865,N159,N1182);
and U281 (N1866,N158,N1182);
not U282 (N1867,N1326);
not U283 (N1868,N1329);
not U284 (N1869,N1332);
not U285 (N1870,N1335);
not U286 (N1871,N1338);
not U287 (N1872,N1341);
not U288 (N1873,N1344);
not U289 (N1874,N1347);
not U290 (N1875,N1350);
not U291 (N1876,N1353);
not U292 (N1877,N1356);
not U293 (N1878,N1359);
not U294 (N1879,N1362);
not U295 (N1880,N1365);
not U296 (N1881,N1368);
not U297 (N1882,N1371);
not U298 (N1883,N1374);
not U299 (N1884,N1377);
buff U300 (N1885,N1199);
buff U301 (N1892,N1194);
buff U302 (N1899,N1199);
buff U303 (N1906,N1194);
not U304 (N1913,N1211);
buff U305 (N1919,N1194);
and U306 (N1926,N44,N1211);
and U307 (N1927,N41,N1211);
and U308 (N1928,N29,N1211);
and U309 (N1929,N26,N1211);
and U310 (N1930,N23,N1211);
not U311 (N1931,N1380);
not U312 (N1932,N1383);
not U313 (N1933,N1386);
not U314 (N1934,N1389);
not U315 (N1935,N1392);
not U316 (N1936,N1395);
not U317 (N1937,N1398);
not U318 (N1938,N1401);
not U319 (N1939,N1404);
not U320 (N1940,N1407);
not U321 (N1941,N1410);
not U322 (N1942,N1413);
not U323 (N1943,N1416);
not U324 (N1944,N1419);
not U325 (N1945,N1422);
not U326 (N1946,N1425);
not U327 (N1947,N1233);
not U328 (N1953,N1244);
and U329 (N1957,N209,N1233);
and U330 (N1958,N216,N1233);
and U331 (N1959,N215,N1233);
and U332 (N1960,N214,N1233);
and U333 (N1961,N213,N1244);
and U334 (N1962,N212,N1244);
and U335 (N1963,N211,N1244);
not U336 (N1965,N1428);
and U337 (N1966,N1222,N636);
not U338 (N1967,N1431);
not U339 (N1968,N1434);
not U340 (N1969,N1437);
not U341 (N1970,N1440);
not U342 (N1971,N1443);
not U343 (N1972,N1446);
not U344 (N1973,N1449);
not U345 (N1974,N1452);
not U346 (N1975,N1455);
not U347 (N1976,N1458);
not U348 (N1977,N1249);
not U349 (N1983,N1256);
and U350 (N1989,N642,N1249);
and U351 (N1990,N644,N1249);
and U352 (N1991,N651,N1249);
and U353 (N1992,N674,N1249);
and U354 (N1993,N660,N1249);
and U355 (N1994,N666,N1256);
and U356 (N1995,N672,N1256);
and U357 (N1996,N673,N1256);
not U358 (N1997,N1263);
buff U359 (N2003,N1194);
and U360 (N2010,N47,N1263);
and U361 (N2011,N35,N1263);
and U362 (N2012,N32,N1263);
and U363 (N2013,N50,N1263);
and U364 (N2014,N66,N1263);
not U365 (N2015,N1461);
not U366 (N2016,N1464);
not U367 (N2017,N1467);
not U368 (N2018,N1470);
not U369 (N2019,N1473);
not U370 (N2020,N1476);
not U371 (N2021,N1479);
not U372 (N2022,N1482);
not U373 (N2023,N1485);
buff U374 (N2024,N1206);
buff U375 (N2031,N1206);
buff U376 (N2038,N1206);
buff U377 (N2045,N1206);
not U378 (N2052,N1270);
not U379 (N2058,N1277);
and U380 (N2064,N706,N1270);
and U381 (N2065,N708,N1270);
and U382 (N2066,N715,N1270);
and U383 (N2067,N721,N1270);
and U384 (N2068,N727,N1270);
and U385 (N2069,N733,N1277);
and U386 (N2070,N734,N1277);
and U387 (N2071,N742,N1277);
and U388 (N2072,N748,N1277);
and U389 (N2073,N749,N1277);
buff U390 (N2074,N1189);
buff U391 (N2081,N1189);
buff U392 (N2086,N1222);
nand U393 (N2107,N1287,N1821);
nand U394 (N2108,N1284,N1822);
not U395 (N2110,N1703);
nand U396 (N2111,N1703,N1832);
nand U397 (N2112,N1308,N1834);
nand U398 (N2113,N1305,N1835);
not U399 (N2114,N1713);
nand U400 (N2115,N1713,N1839);
not U401 (N2117,N1721);
not U402 (N2171,N1758);
nand U403 (N2172,N1758,N1965);
not U404 (N2230,N1708);
buff U405 (N2231,N1537);
buff U406 (N2235,N1551);
or U407 (N2239,N1783,N1782);
or U408 (N2240,N1783,N1125);
or U409 (N2241,N1783,N1793);
or U410 (N2242,N1783,N1794);
or U411 (N2243,N1783,N1795);
or U412 (N2244,N1789,N1796);
or U413 (N2245,N1789,N1797);
or U414 (N2246,N1789,N1798);
or U415 (N2247,N1799,N1811);
or U416 (N2248,N1799,N1812);
or U417 (N2249,N1799,N1813);
or U418 (N2250,N1799,N1814);
or U419 (N2251,N1799,N1815);
or U420 (N2252,N1805,N1816);
or U421 (N2253,N1805,N1817);
or U422 (N2254,N1805,N1818);
or U423 (N2255,N1805,N1819);
or U424 (N2256,N1805,N1820);
nand U425 (N2257,N2107,N2108);
not U426 (N2267,N2074);
nand U427 (N2268,N1299,N2110);
nand U428 (N2269,N2112,N2113);
nand U429 (N2274,N1311,N2114);
not U430 (N2275,N2081);
and U431 (N2277,N141,N1845);
and U432 (N2278,N147,N1845);
and U433 (N2279,N138,N1845);
and U434 (N2280,N144,N1845);
and U435 (N2281,N135,N1845);
and U436 (N2282,N141,N1851);
and U437 (N2283,N147,N1851);
and U438 (N2284,N138,N1851);
and U439 (N2285,N144,N1851);
and U440 (N2286,N135,N1851);
not U441 (N2287,N1885);
not U442 (N2293,N1892);
and U443 (N2299,N103,N1885);
and U444 (N2300,N130,N1885);
and U445 (N2301,N127,N1885);
and U446 (N2302,N124,N1885);
and U447 (N2303,N100,N1885);
and U448 (N2304,N103,N1892);
and U449 (N2305,N130,N1892);
and U450 (N2306,N127,N1892);
and U451 (N2307,N124,N1892);
and U452 (N2308,N100,N1892);
not U453 (N2309,N1899);
not U454 (N2315,N1906);
and U455 (N2321,N115,N1899);
and U456 (N2322,N118,N1899);
and U457 (N2323,N97,N1899);
and U458 (N2324,N94,N1899);
and U459 (N2325,N121,N1899);
and U460 (N2326,N115,N1906);
and U461 (N2327,N118,N1906);
and U462 (N2328,N97,N1906);
and U463 (N2329,N94,N1906);
and U464 (N2330,N121,N1906);
not U465 (N2331,N1919);
and U466 (N2337,N208,N1913);
and U467 (N2338,N198,N1913);
and U468 (N2339,N207,N1913);
and U469 (N2340,N206,N1913);
and U470 (N2341,N205,N1913);
and U471 (N2342,N44,N1919);
and U472 (N2343,N41,N1919);
and U473 (N2344,N29,N1919);
and U474 (N2345,N26,N1919);
and U475 (N2346,N23,N1919);
or U476 (N2347,N1947,N1233);
or U477 (N2348,N1947,N1957);
or U478 (N2349,N1947,N1958);
or U479 (N2350,N1947,N1959);
or U480 (N2351,N1947,N1960);
or U481 (N2352,N1953,N1961);
or U482 (N2353,N1953,N1962);
or U483 (N2354,N1953,N1963);
nand U484 (N2355,N1428,N2171);
not U485 (N2356,N2086);
nand U486 (N2357,N2086,N1967);
and U487 (N2358,N114,N1977);
and U488 (N2359,N113,N1977);
and U489 (N2360,N111,N1977);
and U490 (N2361,N87,N1977);
and U491 (N2362,N112,N1977);
and U492 (N2363,N88,N1983);
and U493 (N2364,N245,N1983);
and U494 (N2365,N271,N1983);
and U495 (N2366,N759,N1983);
and U496 (N2367,N70,N1983);
not U497 (N2368,N2003);
and U498 (N2374,N193,N1997);
and U499 (N2375,N192,N1997);
and U500 (N2376,N191,N1997);
and U501 (N2377,N190,N1997);
and U502 (N2378,N189,N1997);
and U503 (N2379,N47,N2003);
and U504 (N2380,N35,N2003);
and U505 (N2381,N32,N2003);
and U506 (N2382,N50,N2003);
and U507 (N2383,N66,N2003);
not U508 (N2384,N2024);
not U509 (N2390,N2031);
and U510 (N2396,N58,N2024);
and U511 (N2397,N77,N2024);
and U512 (N2398,N78,N2024);
and U513 (N2399,N59,N2024);
and U514 (N2400,N81,N2024);
and U515 (N2401,N80,N2031);
and U516 (N2402,N79,N2031);
and U517 (N2403,N60,N2031);
and U518 (N2404,N61,N2031);
and U519 (N2405,N62,N2031);
not U520 (N2406,N2038);
not U521 (N2412,N2045);
and U522 (N2418,N69,N2038);
and U523 (N2419,N70,N2038);
and U524 (N2420,N74,N2038);
and U525 (N2421,N76,N2038);
and U526 (N2422,N75,N2038);
and U527 (N2423,N73,N2045);
and U528 (N2424,N53,N2045);
and U529 (N2425,N54,N2045);
and U530 (N2426,N55,N2045);
and U531 (N2427,N56,N2045);
and U532 (N2428,N82,N2052);
and U533 (N2429,N65,N2052);
and U534 (N2430,N83,N2052);
and U535 (N2431,N84,N2052);
and U536 (N2432,N85,N2052);
and U537 (N2433,N64,N2058);
and U538 (N2434,N63,N2058);
and U539 (N2435,N86,N2058);
and U540 (N2436,N109,N2058);
and U541 (N2437,N110,N2058);
and U542 (N2441,N2239,N1119);
and U543 (N2442,N2240,N1119);
and U544 (N2446,N2241,N1119);
and U545 (N2450,N2242,N1119);
and U546 (N2454,N2243,N1119);
and U547 (N2458,N2244,N1132);
and U548 (N2462,N2247,N1141);
and U549 (N2466,N2248,N1141);
and U550 (N2470,N2249,N1141);
and U551 (N2474,N2250,N1141);
and U552 (N2478,N2251,N1141);
and U553 (N2482,N2252,N1154);
and U554 (N2488,N2253,N1154);
and U555 (N2496,N2254,N1154);
and U556 (N2502,N2255,N1154);
and U557 (N2508,N2256,N1154);
nand U558 (N2523,N2268,N2111);
nand U559 (N2533,N2274,N2115);
not U560 (N2537,N2235);
or U561 (N2538,N2278,N1858);
or U562 (N2542,N2279,N1859);
or U563 (N2546,N2280,N1860);
or U564 (N2550,N2281,N1861);
or U565 (N2554,N2283,N1863);
or U566 (N2561,N2284,N1864);
or U567 (N2567,N2285,N1865);
or U568 (N2573,N2286,N1866);
or U569 (N2604,N2338,N1927);
or U570 (N2607,N2339,N1928);
or U571 (N2611,N2340,N1929);
or U572 (N2615,N2341,N1930);
and U573 (N2619,N2348,N1227);
and U574 (N2626,N2349,N1227);
and U575 (N2632,N2350,N1227);
and U576 (N2638,N2351,N1227);
and U577 (N2644,N2352,N1240);
nand U578 (N2650,N2355,N2172);
nand U579 (N2653,N1431,N2356);
or U580 (N2654,N2359,N1990);
or U581 (N2658,N2360,N1991);
or U582 (N2662,N2361,N1992);
or U583 (N2666,N2362,N1993);
or U584 (N2670,N2363,N1994);
or U585 (N2674,N2366,N1256);
or U586 (N2680,N2367,N1256);
or U587 (N2688,N2374,N2010);
or U588 (N2692,N2375,N2011);
or U589 (N2696,N2376,N2012);
or U590 (N2700,N2377,N2013);
or U591 (N2704,N2378,N2014);
and U592 (N2728,N2347,N1227);
or U593 (N2729,N2429,N2065);
or U594 (N2733,N2430,N2066);
or U595 (N2737,N2431,N2067);
or U596 (N2741,N2432,N2068);
or U597 (N2745,N2433,N2069);
or U598 (N2749,N2434,N2070);
or U599 (N2753,N2435,N2071);
or U600 (N2757,N2436,N2072);
or U601 (N2761,N2437,N2073);
not U602 (N2765,N2231);
and U603 (N2766,N2354,N1240);
and U604 (N2769,N2353,N1240);
and U605 (N2772,N2246,N1132);
and U606 (N2775,N2245,N1132);
or U607 (N2778,N2282,N1862);
or U608 (N2781,N2358,N1989);
or U609 (N2784,N2365,N1996);
or U610 (N2787,N2364,N1995);
or U611 (N2790,N2337,N1926);
or U612 (N2793,N2277,N1857);
or U613 (N2796,N2428,N2064);
and U614 (N2866,N2257,N1537);
and U615 (N2867,N2257,N1537);
and U616 (N2868,N2257,N1537);
and U617 (N2869,N2257,N1537);
and U618 (N2878,N2269,N1551);
and U619 (N2913,N204,N2287);
and U620 (N2914,N203,N2287);
and U621 (N2915,N202,N2287);
and U622 (N2916,N201,N2287);
and U623 (N2917,N200,N2287);
and U624 (N2918,N235,N2293);
and U625 (N2919,N234,N2293);
and U626 (N2920,N233,N2293);
and U627 (N2921,N232,N2293);
and U628 (N2922,N231,N2293);
and U629 (N2923,N197,N2309);
and U630 (N2924,N187,N2309);
and U631 (N2925,N196,N2309);
and U632 (N2926,N195,N2309);
and U633 (N2927,N194,N2309);
and U634 (N2928,N227,N2315);
and U635 (N2929,N217,N2315);
and U636 (N2930,N226,N2315);
and U637 (N2931,N225,N2315);
and U638 (N2932,N224,N2315);
and U639 (N2933,N239,N2331);
and U640 (N2934,N229,N2331);
and U641 (N2935,N238,N2331);
and U642 (N2936,N237,N2331);
and U643 (N2937,N236,N2331);
nand U644 (N2988,N2653,N2357);
and U645 (N3005,N223,N2368);
and U646 (N3006,N222,N2368);
and U647 (N3007,N221,N2368);
and U648 (N3008,N220,N2368);
and U649 (N3009,N219,N2368);
and U650 (N3020,N812,N2384);
and U651 (N3021,N814,N2384);
and U652 (N3022,N821,N2384);
and U653 (N3023,N827,N2384);
and U654 (N3024,N833,N2384);
and U655 (N3025,N839,N2390);
and U656 (N3026,N845,N2390);
and U657 (N3027,N853,N2390);
and U658 (N3028,N859,N2390);
and U659 (N3029,N865,N2390);
and U660 (N3032,N758,N2406);
and U661 (N3033,N759,N2406);
and U662 (N3034,N762,N2406);
and U663 (N3035,N768,N2406);
and U664 (N3036,N774,N2406);
and U665 (N3037,N780,N2412);
and U666 (N3038,N786,N2412);
and U667 (N3039,N794,N2412);
and U668 (N3040,N800,N2412);
and U669 (N3041,N806,N2412);
buff U670 (N3061,N2257);
buff U671 (N3064,N2257);
buff U672 (N3067,N2269);
buff U673 (N3070,N2269);
not U674 (N3073,N2728);
not U675 (N3080,N2441);
and U676 (N3096,N666,N2644);
and U677 (N3097,N660,N2638);
and U678 (N3101,N1189,N2632);
and U679 (N3107,N651,N2626);
and U680 (N3114,N644,N2619);
and U681 (N3122,N2523,N2257);
or U682 (N3126,N1167,N2866);
and U683 (N3130,N2523,N2257);
or U684 (N3131,N1167,N2869);
and U685 (N3134,N2523,N2257);
not U686 (N3135,N2533);
and U687 (N3136,N666,N2644);
and U688 (N3137,N660,N2638);
and U689 (N3140,N1189,N2632);
and U690 (N3144,N651,N2626);
and U691 (N3149,N644,N2619);
and U692 (N3155,N2533,N2269);
or U693 (N3159,N1174,N2878);
not U694 (N3167,N2778);
and U695 (N3168,N609,N2508);
and U696 (N3169,N604,N2502);
and U697 (N3173,N742,N2496);
and U698 (N3178,N734,N2488);
and U699 (N3184,N599,N2482);
and U700 (N3185,N727,N2573);
and U701 (N3189,N721,N2567);
and U702 (N3195,N715,N2561);
and U703 (N3202,N708,N2554);
and U704 (N3210,N609,N2508);
and U705 (N3211,N604,N2502);
and U706 (N3215,N742,N2496);
and U707 (N3221,N2488,N734);
and U708 (N3228,N599,N2482);
and U709 (N3229,N727,N2573);
and U710 (N3232,N721,N2567);
and U711 (N3236,N715,N2561);
and U712 (N3241,N708,N2554);
or U713 (N3247,N2913,N2299);
or U714 (N3251,N2914,N2300);
or U715 (N3255,N2915,N2301);
or U716 (N3259,N2916,N2302);
or U717 (N3263,N2917,N2303);
or U718 (N3267,N2918,N2304);
or U719 (N3273,N2919,N2305);
or U720 (N3281,N2920,N2306);
or U721 (N3287,N2921,N2307);
or U722 (N3293,N2922,N2308);
or U723 (N3299,N2924,N2322);
or U724 (N3303,N2925,N2323);
or U725 (N3307,N2926,N2324);
or U726 (N3311,N2927,N2325);
or U727 (N3315,N2929,N2327);
or U728 (N3322,N2930,N2328);
or U729 (N3328,N2931,N2329);
or U730 (N3334,N2932,N2330);
or U731 (N3340,N2934,N2343);
or U732 (N3343,N2935,N2344);
or U733 (N3349,N2936,N2345);
or U734 (N3355,N2937,N2346);
and U735 (N3361,N2761,N2478);
and U736 (N3362,N2757,N2474);
and U737 (N3363,N2753,N2470);
and U738 (N3364,N2749,N2466);
and U739 (N3365,N2745,N2462);
and U740 (N3366,N2741,N2550);
and U741 (N3367,N2737,N2546);
and U742 (N3368,N2733,N2542);
and U743 (N3369,N2729,N2538);
and U744 (N3370,N2670,N2458);
and U745 (N3371,N2666,N2454);
and U746 (N3372,N2662,N2450);
and U747 (N3373,N2658,N2446);
and U748 (N3374,N2654,N2442);
and U749 (N3375,N2988,N2650);
and U750 (N3379,N2650,N1966);
not U751 (N3380,N2781);
and U752 (N3381,N695,N2604);
or U753 (N3384,N3005,N2379);
or U754 (N3390,N3006,N2380);
or U755 (N3398,N3007,N2381);
or U756 (N3404,N3008,N2382);
or U757 (N3410,N3009,N2383);
or U758 (N3416,N3021,N2397);
or U759 (N3420,N3022,N2398);
or U760 (N3424,N3023,N2399);
or U761 (N3428,N3024,N2400);
or U762 (N3432,N3025,N2401);
or U763 (N3436,N3026,N2402);
or U764 (N3440,N3027,N2403);
or U765 (N3444,N3028,N2404);
or U766 (N3448,N3029,N2405);
not U767 (N3452,N2790);
not U768 (N3453,N2793);
or U769 (N3454,N3034,N2420);
or U770 (N3458,N3035,N2421);
or U771 (N3462,N3036,N2422);
or U772 (N3466,N3037,N2423);
or U773 (N3470,N3038,N2424);
or U774 (N3474,N3039,N2425);
or U775 (N3478,N3040,N2426);
or U776 (N3482,N3041,N2427);
not U777 (N3486,N2796);
buff U778 (N3487,N2644);
buff U779 (N3490,N2638);
buff U780 (N3493,N2632);
buff U781 (N3496,N2626);
buff U782 (N3499,N2619);
buff U783 (N3502,N2523);
nor U784 (N3507,N1167,N2868);
buff U785 (N3510,N2523);
nor U786 (N3515,N644,N2619);
buff U787 (N3518,N2644);
buff U788 (N3521,N2638);
buff U789 (N3524,N2632);
buff U790 (N3527,N2626);
buff U791 (N3530,N2619);
buff U792 (N3535,N2619);
buff U793 (N3539,N2632);
buff U794 (N3542,N2626);
buff U795 (N3545,N2644);
buff U796 (N3548,N2638);
not U797 (N3551,N2766);
not U798 (N3552,N2769);
buff U799 (N3553,N2442);
buff U800 (N3557,N2450);
buff U801 (N3560,N2446);
buff U802 (N3563,N2458);
buff U803 (N3566,N2454);
not U804 (N3569,N2772);
not U805 (N3570,N2775);
buff U806 (N3571,N2554);
buff U807 (N3574,N2567);
buff U808 (N3577,N2561);
buff U809 (N3580,N2482);
buff U810 (N3583,N2573);
buff U811 (N3586,N2496);
buff U812 (N3589,N2488);
buff U813 (N3592,N2508);
buff U814 (N3595,N2502);
buff U815 (N3598,N2508);
buff U816 (N3601,N2502);
buff U817 (N3604,N2496);
buff U818 (N3607,N2482);
buff U819 (N3610,N2573);
buff U820 (N3613,N2567);
buff U821 (N3616,N2561);
buff U822 (N3619,N2488);
buff U823 (N3622,N2554);
nor U824 (N3625,N734,N2488);
nor U825 (N3628,N708,N2554);
buff U826 (N3631,N2508);
buff U827 (N3634,N2502);
buff U828 (N3637,N2496);
buff U829 (N3640,N2488);
buff U830 (N3643,N2482);
buff U831 (N3646,N2573);
buff U832 (N3649,N2567);
buff U833 (N3652,N2561);
buff U834 (N3655,N2554);
nor U835 (N3658,N2488,N734);
buff U836 (N3661,N2674);
buff U837 (N3664,N2674);
buff U838 (N3667,N2761);
buff U839 (N3670,N2478);
buff U840 (N3673,N2757);
buff U841 (N3676,N2474);
buff U842 (N3679,N2753);
buff U843 (N3682,N2470);
buff U844 (N3685,N2745);
buff U845 (N3688,N2462);
buff U846 (N3691,N2741);
buff U847 (N3694,N2550);
buff U848 (N3697,N2737);
buff U849 (N3700,N2546);
buff U850 (N3703,N2733);
buff U851 (N3706,N2542);
buff U852 (N3709,N2749);
buff U853 (N3712,N2466);
buff U854 (N3715,N2729);
buff U855 (N3718,N2538);
buff U856 (N3721,N2704);
buff U857 (N3724,N2700);
buff U858 (N3727,N2696);
buff U859 (N3730,N2688);
buff U860 (N3733,N2692);
buff U861 (N3736,N2670);
buff U862 (N3739,N2458);
buff U863 (N3742,N2666);
buff U864 (N3745,N2454);
buff U865 (N3748,N2662);
buff U866 (N3751,N2450);
buff U867 (N3754,N2658);
buff U868 (N3757,N2446);
buff U869 (N3760,N2654);
buff U870 (N3763,N2442);
buff U871 (N3766,N2654);
buff U872 (N3769,N2662);
buff U873 (N3772,N2658);
buff U874 (N3775,N2670);
buff U875 (N3778,N2666);
not U876 (N3781,N2784);
not U877 (N3782,N2787);
or U878 (N3783,N2928,N2326);
or U879 (N3786,N2933,N2342);
or U880 (N3789,N2923,N2321);
buff U881 (N3792,N2688);
buff U882 (N3795,N2696);
buff U883 (N3798,N2692);
buff U884 (N3801,N2704);
buff U885 (N3804,N2700);
buff U886 (N3807,N2604);
buff U887 (N3810,N2611);
buff U888 (N3813,N2607);
buff U889 (N3816,N2615);
buff U890 (N3819,N2538);
buff U891 (N3822,N2546);
buff U892 (N3825,N2542);
buff U893 (N3828,N2462);
buff U894 (N3831,N2550);
buff U895 (N3834,N2470);
buff U896 (N3837,N2466);
buff U897 (N3840,N2478);
buff U898 (N3843,N2474);
buff U899 (N3846,N2615);
buff U900 (N3849,N2611);
buff U901 (N3852,N2607);
buff U902 (N3855,N2680);
buff U903 (N3858,N2729);
buff U904 (N3861,N2737);
buff U905 (N3864,N2733);
buff U906 (N3867,N2745);
buff U907 (N3870,N2741);
buff U908 (N3873,N2753);
buff U909 (N3876,N2749);
buff U910 (N3879,N2761);
buff U911 (N3882,N2757);
or U912 (N3885,N3033,N2419);
or U913 (N3888,N3032,N2418);
or U914 (N3891,N3020,N2396);
nand U915 (N3953,N3067,N2117);
not U916 (N3954,N3067);
nand U917 (N3955,N3070,N2537);
not U918 (N3956,N3070);
not U919 (N3958,N3073);
not U920 (N3964,N3080);
or U921 (N4193,N1649,N3379);
or U922 (N4303,N1167,N2867,N3130);
not U923 (N4308,N3061);
not U924 (N4313,N3064);
nand U925 (N4326,N2769,N3551);
nand U926 (N4327,N2766,N3552);
nand U927 (N4333,N2775,N3569);
nand U928 (N4334,N2772,N3570);
nand U929 (N4411,N2787,N3781);
nand U930 (N4412,N2784,N3782);
nand U931 (N4463,N3487,N1828);
not U932 (N4464,N3487);
nand U933 (N4465,N3490,N1829);
not U934 (N4466,N3490);
nand U935 (N4467,N3493,N2267);
not U936 (N4468,N3493);
nand U937 (N4469,N3496,N1830);
not U938 (N4470,N3496);
nand U939 (N4471,N3499,N1833);
not U940 (N4472,N3499);
not U941 (N4473,N3122);
not U942 (N4474,N3126);
nand U943 (N4475,N3518,N1840);
not U944 (N4476,N3518);
nand U945 (N4477,N3521,N1841);
not U946 (N4478,N3521);
nand U947 (N4479,N3524,N2275);
not U948 (N4480,N3524);
nand U949 (N4481,N3527,N1842);
not U950 (N4482,N3527);
nand U951 (N4483,N3530,N1843);
not U952 (N4484,N3530);
not U953 (N4485,N3155);
not U954 (N4486,N3159);
nand U955 (N4487,N1721,N3954);
nand U956 (N4488,N2235,N3956);
not U957 (N4489,N3535);
nand U958 (N4490,N3535,N3958);
not U959 (N4491,N3539);
not U960 (N4492,N3542);
not U961 (N4493,N3545);
not U962 (N4494,N3548);
not U963 (N4495,N3553);
nand U964 (N4496,N3553,N3964);
not U965 (N4497,N3557);
not U966 (N4498,N3560);
not U967 (N4499,N3563);
not U968 (N4500,N3566);
not U969 (N4501,N3571);
nand U970 (N4502,N3571,N3167);
not U971 (N4503,N3574);
not U972 (N4504,N3577);
not U973 (N4505,N3580);
not U974 (N4506,N3583);
nand U975 (N4507,N3598,N1867);
not U976 (N4508,N3598);
nand U977 (N4509,N3601,N1868);
not U978 (N4510,N3601);
nand U979 (N4511,N3604,N1869);
not U980 (N4512,N3604);
nand U981 (N4513,N3607,N1870);
not U982 (N4514,N3607);
nand U983 (N4515,N3610,N1871);
not U984 (N4516,N3610);
nand U985 (N4517,N3613,N1872);
not U986 (N4518,N3613);
nand U987 (N4519,N3616,N1873);
not U988 (N4520,N3616);
nand U989 (N4521,N3619,N1874);
not U990 (N4522,N3619);
nand U991 (N4523,N3622,N1875);
not U992 (N4524,N3622);
nand U993 (N4525,N3631,N1876);
not U994 (N4526,N3631);
nand U995 (N4527,N3634,N1877);
not U996 (N4528,N3634);
nand U997 (N4529,N3637,N1878);
not U998 (N4530,N3637);
nand U999 (N4531,N3640,N1879);
not U1000 (N4532,N3640);
nand U1001 (N4533,N3643,N1880);
not U1002 (N4534,N3643);
nand U1003 (N4535,N3646,N1881);
not U1004 (N4536,N3646);
nand U1005 (N4537,N3649,N1882);
not U1006 (N4538,N3649);
nand U1007 (N4539,N3652,N1883);
not U1008 (N4540,N3652);
nand U1009 (N4541,N3655,N1884);
not U1010 (N4542,N3655);
not U1011 (N4543,N3658);
and U1012 (N4544,N806,N3293);
and U1013 (N4545,N800,N3287);
and U1014 (N4549,N794,N3281);
and U1015 (N4555,N3273,N786);
and U1016 (N4562,N780,N3267);
and U1017 (N4563,N774,N3355);
and U1018 (N4566,N768,N3349);
and U1019 (N4570,N762,N3343);
not U1020 (N4575,N3661);
and U1021 (N4576,N806,N3293);
and U1022 (N4577,N800,N3287);
and U1023 (N4581,N794,N3281);
and U1024 (N4586,N786,N3273);
and U1025 (N4592,N780,N3267);
and U1026 (N4593,N774,N3355);
and U1027 (N4597,N768,N3349);
and U1028 (N4603,N762,N3343);
not U1029 (N4610,N3664);
not U1030 (N4611,N3667);
not U1031 (N4612,N3670);
not U1032 (N4613,N3673);
not U1033 (N4614,N3676);
not U1034 (N4615,N3679);
not U1035 (N4616,N3682);
not U1036 (N4617,N3685);
not U1037 (N4618,N3688);
not U1038 (N4619,N3691);
not U1039 (N4620,N3694);
not U1040 (N4621,N3697);
not U1041 (N4622,N3700);
not U1042 (N4623,N3703);
not U1043 (N4624,N3706);
not U1044 (N4625,N3709);
not U1045 (N4626,N3712);
not U1046 (N4627,N3715);
not U1047 (N4628,N3718);
not U1048 (N4629,N3721);
and U1049 (N4630,N3448,N2704);
not U1050 (N4631,N3724);
and U1051 (N4632,N3444,N2700);
not U1052 (N4633,N3727);
and U1053 (N4634,N3440,N2696);
and U1054 (N4635,N3436,N2692);
not U1055 (N4636,N3730);
and U1056 (N4637,N3432,N2688);
and U1057 (N4638,N3428,N3311);
and U1058 (N4639,N3424,N3307);
and U1059 (N4640,N3420,N3303);
and U1060 (N4641,N3416,N3299);
not U1061 (N4642,N3733);
not U1062 (N4643,N3736);
not U1063 (N4644,N3739);
not U1064 (N4645,N3742);
not U1065 (N4646,N3745);
not U1066 (N4647,N3748);
not U1067 (N4648,N3751);
not U1068 (N4649,N3754);
not U1069 (N4650,N3757);
not U1070 (N4651,N3760);
not U1071 (N4652,N3763);
not U1072 (N4653,N3375);
and U1073 (N4656,N865,N3410);
and U1074 (N4657,N859,N3404);
and U1075 (N4661,N853,N3398);
and U1076 (N4667,N3390,N845);
and U1077 (N4674,N839,N3384);
and U1078 (N4675,N833,N3334);
and U1079 (N4678,N827,N3328);
and U1080 (N4682,N821,N3322);
and U1081 (N4687,N814,N3315);
not U1082 (N4693,N3766);
nand U1083 (N4694,N3766,N3380);
not U1084 (N4695,N3769);
not U1085 (N4696,N3772);
not U1086 (N4697,N3775);
not U1087 (N4698,N3778);
not U1088 (N4699,N3783);
not U1089 (N4700,N3786);
and U1090 (N4701,N865,N3410);
and U1091 (N4702,N859,N3404);
and U1092 (N4706,N853,N3398);
and U1093 (N4711,N845,N3390);
and U1094 (N4717,N839,N3384);
and U1095 (N4718,N833,N3334);
and U1096 (N4722,N827,N3328);
and U1097 (N4728,N821,N3322);
and U1098 (N4735,N814,N3315);
not U1099 (N4743,N3789);
not U1100 (N4744,N3792);
not U1101 (N4745,N3807);
nand U1102 (N4746,N3807,N3452);
not U1103 (N4747,N3810);
not U1104 (N4748,N3813);
not U1105 (N4749,N3816);
not U1106 (N4750,N3819);
nand U1107 (N4751,N3819,N3453);
not U1108 (N4752,N3822);
not U1109 (N4753,N3825);
not U1110 (N4754,N3828);
not U1111 (N4755,N3831);
and U1112 (N4756,N3482,N3263);
and U1113 (N4757,N3478,N3259);
and U1114 (N4758,N3474,N3255);
and U1115 (N4759,N3470,N3251);
and U1116 (N4760,N3466,N3247);
not U1117 (N4761,N3846);
and U1118 (N4762,N3462,N2615);
not U1119 (N4763,N3849);
and U1120 (N4764,N3458,N2611);
not U1121 (N4765,N3852);
and U1122 (N4766,N3454,N2607);
and U1123 (N4767,N2680,N3381);
not U1124 (N4768,N3855);
and U1125 (N4769,N3340,N695);
not U1126 (N4775,N3858);
nand U1127 (N4776,N3858,N3486);
not U1128 (N4777,N3861);
not U1129 (N4778,N3864);
not U1130 (N4779,N3867);
not U1131 (N4780,N3870);
not U1132 (N4781,N3885);
not U1133 (N4782,N3888);
not U1134 (N4783,N3891);
or U1135 (N4784,N3131,N3134);
not U1136 (N4789,N3502);
not U1137 (N4790,N3131);
not U1138 (N4793,N3507);
not U1139 (N4794,N3510);
not U1140 (N4795,N3515);
buff U1141 (N4796,N3114);
not U1142 (N4799,N3586);
not U1143 (N4800,N3589);
not U1144 (N4801,N3592);
not U1145 (N4802,N3595);
nand U1146 (N4803,N4326,N4327);
nand U1147 (N4806,N4333,N4334);
not U1148 (N4809,N3625);
buff U1149 (N4810,N3178);
not U1150 (N4813,N3628);
buff U1151 (N4814,N3202);
buff U1152 (N4817,N3221);
buff U1153 (N4820,N3293);
buff U1154 (N4823,N3287);
buff U1155 (N4826,N3281);
buff U1156 (N4829,N3273);
buff U1157 (N4832,N3267);
buff U1158 (N4835,N3355);
buff U1159 (N4838,N3349);
buff U1160 (N4841,N3343);
nor U1161 (N4844,N3273,N786);
buff U1162 (N4847,N3293);
buff U1163 (N4850,N3287);
buff U1164 (N4853,N3281);
buff U1165 (N4856,N3267);
buff U1166 (N4859,N3355);
buff U1167 (N4862,N3349);
buff U1168 (N4865,N3343);
buff U1169 (N4868,N3273);
nor U1170 (N4871,N786,N3273);
buff U1171 (N4874,N3448);
buff U1172 (N4877,N3444);
buff U1173 (N4880,N3440);
buff U1174 (N4883,N3432);
buff U1175 (N4886,N3428);
buff U1176 (N4889,N3311);
buff U1177 (N4892,N3424);
buff U1178 (N4895,N3307);
buff U1179 (N4898,N3420);
buff U1180 (N4901,N3303);
buff U1181 (N4904,N3436);
buff U1182 (N4907,N3416);
buff U1183 (N4910,N3299);
buff U1184 (N4913,N3410);
buff U1185 (N4916,N3404);
buff U1186 (N4919,N3398);
buff U1187 (N4922,N3390);
buff U1188 (N4925,N3384);
buff U1189 (N4928,N3334);
buff U1190 (N4931,N3328);
buff U1191 (N4934,N3322);
buff U1192 (N4937,N3315);
nor U1193 (N4940,N3390,N845);
buff U1194 (N4943,N3315);
buff U1195 (N4946,N3328);
buff U1196 (N4949,N3322);
buff U1197 (N4952,N3384);
buff U1198 (N4955,N3334);
buff U1199 (N4958,N3398);
buff U1200 (N4961,N3390);
buff U1201 (N4964,N3410);
buff U1202 (N4967,N3404);
buff U1203 (N4970,N3340);
buff U1204 (N4973,N3349);
buff U1205 (N4976,N3343);
buff U1206 (N4979,N3267);
buff U1207 (N4982,N3355);
buff U1208 (N4985,N3281);
buff U1209 (N4988,N3273);
buff U1210 (N4991,N3293);
buff U1211 (N4994,N3287);
nand U1212 (N4997,N4411,N4412);
buff U1213 (N5000,N3410);
buff U1214 (N5003,N3404);
buff U1215 (N5006,N3398);
buff U1216 (N5009,N3384);
buff U1217 (N5012,N3334);
buff U1218 (N5015,N3328);
buff U1219 (N5018,N3322);
buff U1220 (N5021,N3390);
buff U1221 (N5024,N3315);
nor U1222 (N5027,N845,N3390);
nor U1223 (N5030,N814,N3315);
buff U1224 (N5033,N3299);
buff U1225 (N5036,N3307);
buff U1226 (N5039,N3303);
buff U1227 (N5042,N3311);
not U1228 (N5045,N3795);
not U1229 (N5046,N3798);
not U1230 (N5047,N3801);
not U1231 (N5048,N3804);
buff U1232 (N5049,N3247);
buff U1233 (N5052,N3255);
buff U1234 (N5055,N3251);
buff U1235 (N5058,N3263);
buff U1236 (N5061,N3259);
not U1237 (N5064,N3834);
not U1238 (N5065,N3837);
not U1239 (N5066,N3840);
not U1240 (N5067,N3843);
buff U1241 (N5068,N3482);
buff U1242 (N5071,N3263);
buff U1243 (N5074,N3478);
buff U1244 (N5077,N3259);
buff U1245 (N5080,N3474);
buff U1246 (N5083,N3255);
buff U1247 (N5086,N3466);
buff U1248 (N5089,N3247);
buff U1249 (N5092,N3462);
buff U1250 (N5095,N3458);
buff U1251 (N5098,N3454);
buff U1252 (N5101,N3470);
buff U1253 (N5104,N3251);
buff U1254 (N5107,N3381);
not U1255 (N5110,N3873);
not U1256 (N5111,N3876);
not U1257 (N5112,N3879);
not U1258 (N5113,N3882);
buff U1259 (N5114,N3458);
buff U1260 (N5117,N3454);
buff U1261 (N5120,N3466);
buff U1262 (N5123,N3462);
buff U1263 (N5126,N3474);
buff U1264 (N5129,N3470);
buff U1265 (N5132,N3482);
buff U1266 (N5135,N3478);
buff U1267 (N5138,N3416);
buff U1268 (N5141,N3424);
buff U1269 (N5144,N3420);
buff U1270 (N5147,N3432);
buff U1271 (N5150,N3428);
buff U1272 (N5153,N3440);
buff U1273 (N5156,N3436);
buff U1274 (N5159,N3448);
buff U1275 (N5162,N3444);
nand U1276 (N5165,N4486,N4485);
nand U1277 (N5166,N4474,N4473);
nand U1278 (N5167,N1290,N4464);
nand U1279 (N5168,N1293,N4466);
nand U1280 (N5169,N2074,N4468);
nand U1281 (N5170,N1296,N4470);
nand U1282 (N5171,N1302,N4472);
nand U1283 (N5172,N1314,N4476);
nand U1284 (N5173,N1317,N4478);
nand U1285 (N5174,N2081,N4480);
nand U1286 (N5175,N1320,N4482);
nand U1287 (N5176,N1323,N4484);
nand U1288 (N5177,N3953,N4487);
nand U1289 (N5178,N3955,N4488);
nand U1290 (N5179,N3073,N4489);
nand U1291 (N5180,N3542,N4491);
nand U1292 (N5181,N3539,N4492);
nand U1293 (N5182,N3548,N4493);
nand U1294 (N5183,N3545,N4494);
nand U1295 (N5184,N3080,N4495);
nand U1296 (N5185,N3560,N4497);
nand U1297 (N5186,N3557,N4498);
nand U1298 (N5187,N3566,N4499);
nand U1299 (N5188,N3563,N4500);
nand U1300 (N5189,N2778,N4501);
nand U1301 (N5190,N3577,N4503);
nand U1302 (N5191,N3574,N4504);
nand U1303 (N5192,N3583,N4505);
nand U1304 (N5193,N3580,N4506);
nand U1305 (N5196,N1326,N4508);
nand U1306 (N5197,N1329,N4510);
nand U1307 (N5198,N1332,N4512);
nand U1308 (N5199,N1335,N4514);
nand U1309 (N5200,N1338,N4516);
nand U1310 (N5201,N1341,N4518);
nand U1311 (N5202,N1344,N4520);
nand U1312 (N5203,N1347,N4522);
nand U1313 (N5204,N1350,N4524);
nand U1314 (N5205,N1353,N4526);
nand U1315 (N5206,N1356,N4528);
nand U1316 (N5207,N1359,N4530);
nand U1317 (N5208,N1362,N4532);
nand U1318 (N5209,N1365,N4534);
nand U1319 (N5210,N1368,N4536);
nand U1320 (N5211,N1371,N4538);
nand U1321 (N5212,N1374,N4540);
nand U1322 (N5213,N1377,N4542);
nand U1323 (N5283,N3670,N4611);
nand U1324 (N5284,N3667,N4612);
nand U1325 (N5285,N3676,N4613);
nand U1326 (N5286,N3673,N4614);
nand U1327 (N5287,N3682,N4615);
nand U1328 (N5288,N3679,N4616);
nand U1329 (N5289,N3688,N4617);
nand U1330 (N5290,N3685,N4618);
nand U1331 (N5291,N3694,N4619);
nand U1332 (N5292,N3691,N4620);
nand U1333 (N5293,N3700,N4621);
nand U1334 (N5294,N3697,N4622);
nand U1335 (N5295,N3706,N4623);
nand U1336 (N5296,N3703,N4624);
nand U1337 (N5297,N3712,N4625);
nand U1338 (N5298,N3709,N4626);
nand U1339 (N5299,N3718,N4627);
nand U1340 (N5300,N3715,N4628);
nand U1341 (N5314,N3739,N4643);
nand U1342 (N5315,N3736,N4644);
nand U1343 (N5316,N3745,N4645);
nand U1344 (N5317,N3742,N4646);
nand U1345 (N5318,N3751,N4647);
nand U1346 (N5319,N3748,N4648);
nand U1347 (N5320,N3757,N4649);
nand U1348 (N5321,N3754,N4650);
nand U1349 (N5322,N3763,N4651);
nand U1350 (N5323,N3760,N4652);
not U1351 (N5324,N4193);
nand U1352 (N5363,N2781,N4693);
nand U1353 (N5364,N3772,N4695);
nand U1354 (N5365,N3769,N4696);
nand U1355 (N5366,N3778,N4697);
nand U1356 (N5367,N3775,N4698);
nand U1357 (N5425,N2790,N4745);
nand U1358 (N5426,N3813,N4747);
nand U1359 (N5427,N3810,N4748);
nand U1360 (N5429,N2793,N4750);
nand U1361 (N5430,N3825,N4752);
nand U1362 (N5431,N3822,N4753);
nand U1363 (N5432,N3831,N4754);
nand U1364 (N5433,N3828,N4755);
nand U1365 (N5451,N2796,N4775);
nand U1366 (N5452,N3864,N4777);
nand U1367 (N5453,N3861,N4778);
nand U1368 (N5454,N3870,N4779);
nand U1369 (N5455,N3867,N4780);
nand U1370 (N5456,N3888,N4781);
nand U1371 (N5457,N3885,N4782);
not U1372 (N5469,N4303);
nand U1373 (N5474,N3589,N4799);
nand U1374 (N5475,N3586,N4800);
nand U1375 (N5476,N3595,N4801);
nand U1376 (N5477,N3592,N4802);
nand U1377 (N5571,N3798,N5045);
nand U1378 (N5572,N3795,N5046);
nand U1379 (N5573,N3804,N5047);
nand U1380 (N5574,N3801,N5048);
nand U1381 (N5584,N3837,N5064);
nand U1382 (N5585,N3834,N5065);
nand U1383 (N5586,N3843,N5066);
nand U1384 (N5587,N3840,N5067);
nand U1385 (N5602,N3876,N5110);
nand U1386 (N5603,N3873,N5111);
nand U1387 (N5604,N3882,N5112);
nand U1388 (N5605,N3879,N5113);
nand U1389 (N5631,N5324,N4653);
nand U1390 (N5632,N4463,N5167);
nand U1391 (N5640,N4465,N5168);
nand U1392 (N5654,N4467,N5169);
nand U1393 (N5670,N4469,N5170);
nand U1394 (N5683,N4471,N5171);
nand U1395 (N5690,N4475,N5172);
nand U1396 (N5697,N4477,N5173);
nand U1397 (N5707,N4479,N5174);
nand U1398 (N5718,N4481,N5175);
nand U1399 (N5728,N4483,N5176);
not U1400 (N5735,N5177);
nand U1401 (N5736,N5179,N4490);
nand U1402 (N5740,N5180,N5181);
nand U1403 (N5744,N5182,N5183);
nand U1404 (N5747,N5184,N4496);
nand U1405 (N5751,N5185,N5186);
nand U1406 (N5755,N5187,N5188);
nand U1407 (N5758,N5189,N4502);
nand U1408 (N5762,N5190,N5191);
nand U1409 (N5766,N5192,N5193);
not U1410 (N5769,N4803);
not U1411 (N5770,N4806);
nand U1412 (N5771,N4507,N5196);
nand U1413 (N5778,N4509,N5197);
nand U1414 (N5789,N4511,N5198);
nand U1415 (N5799,N4513,N5199);
nand U1416 (N5807,N4515,N5200);
nand U1417 (N5821,N4517,N5201);
nand U1418 (N5837,N4519,N5202);
nand U1419 (N5850,N4521,N5203);
nand U1420 (N5856,N4523,N5204);
nand U1421 (N5863,N4525,N5205);
nand U1422 (N5870,N4527,N5206);
nand U1423 (N5881,N4529,N5207);
nand U1424 (N5892,N4531,N5208);
nand U1425 (N5898,N4533,N5209);
nand U1426 (N5905,N4535,N5210);
nand U1427 (N5915,N4537,N5211);
nand U1428 (N5926,N4539,N5212);
nand U1429 (N5936,N4541,N5213);
not U1430 (N5943,N4817);
nand U1431 (N5944,N4820,N1931);
not U1432 (N5945,N4820);
nand U1433 (N5946,N4823,N1932);
not U1434 (N5947,N4823);
nand U1435 (N5948,N4826,N1933);
not U1436 (N5949,N4826);
nand U1437 (N5950,N4829,N1934);
not U1438 (N5951,N4829);
nand U1439 (N5952,N4832,N1935);
not U1440 (N5953,N4832);
nand U1441 (N5954,N4835,N1936);
not U1442 (N5955,N4835);
nand U1443 (N5956,N4838,N1937);
not U1444 (N5957,N4838);
nand U1445 (N5958,N4841,N1938);
not U1446 (N5959,N4841);
and U1447 (N5960,N2674,N4769);
not U1448 (N5966,N4844);
nand U1449 (N5967,N4847,N1939);
not U1450 (N5968,N4847);
nand U1451 (N5969,N4850,N1940);
not U1452 (N5970,N4850);
nand U1453 (N5971,N4853,N1941);
not U1454 (N5972,N4853);
nand U1455 (N5973,N4856,N1942);
not U1456 (N5974,N4856);
nand U1457 (N5975,N4859,N1943);
not U1458 (N5976,N4859);
nand U1459 (N5977,N4862,N1944);
not U1460 (N5978,N4862);
nand U1461 (N5979,N4865,N1945);
not U1462 (N5980,N4865);
and U1463 (N5981,N2674,N4769);
nand U1464 (N5989,N4868,N1946);
not U1465 (N5990,N4868);
nand U1466 (N5991,N5283,N5284);
nand U1467 (N5996,N5285,N5286);
nand U1468 (N6000,N5287,N5288);
nand U1469 (N6003,N5289,N5290);
nand U1470 (N6009,N5291,N5292);
nand U1471 (N6014,N5293,N5294);
nand U1472 (N6018,N5295,N5296);
nand U1473 (N6021,N5297,N5298);
nand U1474 (N6022,N5299,N5300);
not U1475 (N6023,N4874);
nand U1476 (N6024,N4874,N4629);
not U1477 (N6025,N4877);
nand U1478 (N6026,N4877,N4631);
not U1479 (N6027,N4880);
nand U1480 (N6028,N4880,N4633);
not U1481 (N6029,N4883);
nand U1482 (N6030,N4883,N4636);
not U1483 (N6031,N4886);
not U1484 (N6032,N4889);
not U1485 (N6033,N4892);
not U1486 (N6034,N4895);
not U1487 (N6035,N4898);
not U1488 (N6036,N4901);
not U1489 (N6037,N4904);
nand U1490 (N6038,N4904,N4642);
not U1491 (N6039,N4907);
not U1492 (N6040,N4910);
nand U1493 (N6041,N5314,N5315);
nand U1494 (N6047,N5316,N5317);
nand U1495 (N6052,N5318,N5319);
nand U1496 (N6056,N5320,N5321);
nand U1497 (N6059,N5322,N5323);
nand U1498 (N6060,N4913,N1968);
not U1499 (N6061,N4913);
nand U1500 (N6062,N4916,N1969);
not U1501 (N6063,N4916);
nand U1502 (N6064,N4919,N1970);
not U1503 (N6065,N4919);
nand U1504 (N6066,N4922,N1971);
not U1505 (N6067,N4922);
nand U1506 (N6068,N4925,N1972);
not U1507 (N6069,N4925);
nand U1508 (N6070,N4928,N1973);
not U1509 (N6071,N4928);
nand U1510 (N6072,N4931,N1974);
not U1511 (N6073,N4931);
nand U1512 (N6074,N4934,N1975);
not U1513 (N6075,N4934);
nand U1514 (N6076,N4937,N1976);
not U1515 (N6077,N4937);
not U1516 (N6078,N4940);
nand U1517 (N6079,N5363,N4694);
nand U1518 (N6083,N5364,N5365);
nand U1519 (N6087,N5366,N5367);
not U1520 (N6090,N4943);
nand U1521 (N6091,N4943,N4699);
not U1522 (N6092,N4946);
not U1523 (N6093,N4949);
not U1524 (N6094,N4952);
not U1525 (N6095,N4955);
not U1526 (N6096,N4970);
nand U1527 (N6097,N4970,N4700);
not U1528 (N6098,N4973);
not U1529 (N6099,N4976);
not U1530 (N6100,N4979);
not U1531 (N6101,N4982);
not U1532 (N6102,N4997);
nand U1533 (N6103,N5000,N2015);
not U1534 (N6104,N5000);
nand U1535 (N6105,N5003,N2016);
not U1536 (N6106,N5003);
nand U1537 (N6107,N5006,N2017);
not U1538 (N6108,N5006);
nand U1539 (N6109,N5009,N2018);
not U1540 (N6110,N5009);
nand U1541 (N6111,N5012,N2019);
not U1542 (N6112,N5012);
nand U1543 (N6113,N5015,N2020);
not U1544 (N6114,N5015);
nand U1545 (N6115,N5018,N2021);
not U1546 (N6116,N5018);
nand U1547 (N6117,N5021,N2022);
not U1548 (N6118,N5021);
nand U1549 (N6119,N5024,N2023);
not U1550 (N6120,N5024);
not U1551 (N6121,N5033);
nand U1552 (N6122,N5033,N4743);
not U1553 (N6123,N5036);
not U1554 (N6124,N5039);
nand U1555 (N6125,N5042,N4744);
not U1556 (N6126,N5042);
nand U1557 (N6127,N5425,N4746);
nand U1558 (N6131,N5426,N5427);
not U1559 (N6135,N5049);
nand U1560 (N6136,N5049,N4749);
nand U1561 (N6137,N5429,N4751);
nand U1562 (N6141,N5430,N5431);
nand U1563 (N6145,N5432,N5433);
not U1564 (N6148,N5068);
not U1565 (N6149,N5071);
not U1566 (N6150,N5074);
not U1567 (N6151,N5077);
not U1568 (N6152,N5080);
not U1569 (N6153,N5083);
not U1570 (N6154,N5086);
not U1571 (N6155,N5089);
not U1572 (N6156,N5092);
nand U1573 (N6157,N5092,N4761);
not U1574 (N6158,N5095);
nand U1575 (N6159,N5095,N4763);
not U1576 (N6160,N5098);
nand U1577 (N6161,N5098,N4765);
not U1578 (N6162,N5101);
not U1579 (N6163,N5104);
nand U1580 (N6164,N5107,N4768);
not U1581 (N6165,N5107);
nand U1582 (N6166,N5451,N4776);
nand U1583 (N6170,N5452,N5453);
nand U1584 (N6174,N5454,N5455);
nand U1585 (N6177,N5456,N5457);
not U1586 (N6181,N5114);
not U1587 (N6182,N5117);
not U1588 (N6183,N5120);
not U1589 (N6184,N5123);
not U1590 (N6185,N5138);
nand U1591 (N6186,N5138,N4783);
not U1592 (N6187,N5141);
not U1593 (N6188,N5144);
not U1594 (N6189,N5147);
not U1595 (N6190,N5150);
not U1596 (N6191,N4784);
nand U1597 (N6192,N4784,N2230);
not U1598 (N6193,N4790);
nand U1599 (N6194,N4790,N2765);
not U1600 (N6195,N4796);
nand U1601 (N6196,N5476,N5477);
nand U1602 (N6199,N5474,N5475);
not U1603 (N6202,N4810);
not U1604 (N6203,N4814);
buff U1605 (N6204,N4769);
buff U1606 (N6207,N4555);
buff U1607 (N6210,N4769);
not U1608 (N6213,N4871);
buff U1609 (N6214,N4586);
nor U1610 (N6217,N2674,N4769);
buff U1611 (N6220,N4667);
not U1612 (N6223,N4958);
not U1613 (N6224,N4961);
not U1614 (N6225,N4964);
not U1615 (N6226,N4967);
not U1616 (N6227,N4985);
not U1617 (N6228,N4988);
not U1618 (N6229,N4991);
not U1619 (N6230,N4994);
not U1620 (N6231,N5027);
buff U1621 (N6232,N4711);
not U1622 (N6235,N5030);
buff U1623 (N6236,N4735);
not U1624 (N6239,N5052);
not U1625 (N6240,N5055);
not U1626 (N6241,N5058);
not U1627 (N6242,N5061);
nand U1628 (N6243,N5573,N5574);
nand U1629 (N6246,N5571,N5572);
nand U1630 (N6249,N5586,N5587);
nand U1631 (N6252,N5584,N5585);
not U1632 (N6255,N5126);
not U1633 (N6256,N5129);
not U1634 (N6257,N5132);
not U1635 (N6258,N5135);
not U1636 (N6259,N5153);
not U1637 (N6260,N5156);
not U1638 (N6261,N5159);
not U1639 (N6262,N5162);
nand U1640 (N6263,N5604,N5605);
nand U1641 (N6266,N5602,N5603);
nand U1642 (N6540,N1380,N5945);
nand U1643 (N6541,N1383,N5947);
nand U1644 (N6542,N1386,N5949);
nand U1645 (N6543,N1389,N5951);
nand U1646 (N6544,N1392,N5953);
nand U1647 (N6545,N1395,N5955);
nand U1648 (N6546,N1398,N5957);
nand U1649 (N6547,N1401,N5959);
nand U1650 (N6555,N1404,N5968);
nand U1651 (N6556,N1407,N5970);
nand U1652 (N6557,N1410,N5972);
nand U1653 (N6558,N1413,N5974);
nand U1654 (N6559,N1416,N5976);
nand U1655 (N6560,N1419,N5978);
nand U1656 (N6561,N1422,N5980);
nand U1657 (N6569,N1425,N5990);
nand U1658 (N6594,N3721,N6023);
nand U1659 (N6595,N3724,N6025);
nand U1660 (N6596,N3727,N6027);
nand U1661 (N6597,N3730,N6029);
nand U1662 (N6598,N4889,N6031);
nand U1663 (N6599,N4886,N6032);
nand U1664 (N6600,N4895,N6033);
nand U1665 (N6601,N4892,N6034);
nand U1666 (N6602,N4901,N6035);
nand U1667 (N6603,N4898,N6036);
nand U1668 (N6604,N3733,N6037);
nand U1669 (N6605,N4910,N6039);
nand U1670 (N6606,N4907,N6040);
nand U1671 (N6621,N1434,N6061);
nand U1672 (N6622,N1437,N6063);
nand U1673 (N6623,N1440,N6065);
nand U1674 (N6624,N1443,N6067);
nand U1675 (N6625,N1446,N6069);
nand U1676 (N6626,N1449,N6071);
nand U1677 (N6627,N1452,N6073);
nand U1678 (N6628,N1455,N6075);
nand U1679 (N6629,N1458,N6077);
nand U1680 (N6639,N3783,N6090);
nand U1681 (N6640,N4949,N6092);
nand U1682 (N6641,N4946,N6093);
nand U1683 (N6642,N4955,N6094);
nand U1684 (N6643,N4952,N6095);
nand U1685 (N6644,N3786,N6096);
nand U1686 (N6645,N4976,N6098);
nand U1687 (N6646,N4973,N6099);
nand U1688 (N6647,N4982,N6100);
nand U1689 (N6648,N4979,N6101);
nand U1690 (N6649,N1461,N6104);
nand U1691 (N6650,N1464,N6106);
nand U1692 (N6651,N1467,N6108);
nand U1693 (N6652,N1470,N6110);
nand U1694 (N6653,N1473,N6112);
nand U1695 (N6654,N1476,N6114);
nand U1696 (N6655,N1479,N6116);
nand U1697 (N6656,N1482,N6118);
nand U1698 (N6657,N1485,N6120);
nand U1699 (N6658,N3789,N6121);
nand U1700 (N6659,N5039,N6123);
nand U1701 (N6660,N5036,N6124);
nand U1702 (N6661,N3792,N6126);
nand U1703 (N6668,N3816,N6135);
nand U1704 (N6677,N5071,N6148);
nand U1705 (N6678,N5068,N6149);
nand U1706 (N6679,N5077,N6150);
nand U1707 (N6680,N5074,N6151);
nand U1708 (N6681,N5083,N6152);
nand U1709 (N6682,N5080,N6153);
nand U1710 (N6683,N5089,N6154);
nand U1711 (N6684,N5086,N6155);
nand U1712 (N6685,N3846,N6156);
nand U1713 (N6686,N3849,N6158);
nand U1714 (N6687,N3852,N6160);
nand U1715 (N6688,N5104,N6162);
nand U1716 (N6689,N5101,N6163);
nand U1717 (N6690,N3855,N6165);
nand U1718 (N6702,N5117,N6181);
nand U1719 (N6703,N5114,N6182);
nand U1720 (N6704,N5123,N6183);
nand U1721 (N6705,N5120,N6184);
nand U1722 (N6706,N3891,N6185);
nand U1723 (N6707,N5144,N6187);
nand U1724 (N6708,N5141,N6188);
nand U1725 (N6709,N5150,N6189);
nand U1726 (N6710,N5147,N6190);
nand U1727 (N6711,N1708,N6191);
nand U1728 (N6712,N2231,N6193);
nand U1729 (N6729,N4961,N6223);
nand U1730 (N6730,N4958,N6224);
nand U1731 (N6731,N4967,N6225);
nand U1732 (N6732,N4964,N6226);
nand U1733 (N6733,N4988,N6227);
nand U1734 (N6734,N4985,N6228);
nand U1735 (N6735,N4994,N6229);
nand U1736 (N6736,N4991,N6230);
nand U1737 (N6741,N5055,N6239);
nand U1738 (N6742,N5052,N6240);
nand U1739 (N6743,N5061,N6241);
nand U1740 (N6744,N5058,N6242);
nand U1741 (N6751,N5129,N6255);
nand U1742 (N6752,N5126,N6256);
nand U1743 (N6753,N5135,N6257);
nand U1744 (N6754,N5132,N6258);
nand U1745 (N6755,N5156,N6259);
nand U1746 (N6756,N5153,N6260);
nand U1747 (N6757,N5162,N6261);
nand U1748 (N6758,N5159,N6262);
not U1749 (N6761,N5892);
and U1750 (N6762,N5683,N5670,N5654,N5640,N5632);
and U1751 (N6766,N5632,N3097);
and U1752 (N6767,N5640,N5632,N3101);
and U1753 (N6768,N5654,N5632,N3107,N5640);
and U1754 (N6769,N5670,N5654,N5632,N3114,N5640);
and U1755 (N6770,N5640,N3101);
and U1756 (N6771,N5654,N3107,N5640);
and U1757 (N6772,N5670,N5654,N3114,N5640);
and U1758 (N6773,N5683,N5654,N5640,N5670);
and U1759 (N6774,N5640,N3101);
and U1760 (N6775,N5654,N3107,N5640);
and U1761 (N6776,N5670,N5654,N3114,N5640);
and U1762 (N6777,N5654,N3107);
and U1763 (N6778,N5670,N5654,N3114);
and U1764 (N6779,N5683,N5654,N5670);
and U1765 (N6780,N5654,N3107);
and U1766 (N6781,N5670,N5654,N3114);
and U1767 (N6782,N5670,N3114);
and U1768 (N6783,N5683,N5670);
and U1769 (N6784,N5697,N5728,N5707,N5690,N5718);
and U1770 (N6787,N5690,N3137);
and U1771 (N6788,N5697,N5690,N3140);
and U1772 (N6789,N5707,N5690,N3144,N5697);
and U1773 (N6790,N5718,N5707,N5690,N3149,N5697);
and U1774 (N6791,N5697,N3140);
and U1775 (N6792,N5707,N3144,N5697);
and U1776 (N6793,N5718,N5707,N3149,N5697);
and U1777 (N6794,N3144,N5707);
and U1778 (N6795,N5718,N5707,N3149);
and U1779 (N6796,N5718,N3149);
not U1780 (N6797,N5736);
not U1781 (N6800,N5740);
not U1782 (N6803,N5747);
not U1783 (N6806,N5751);
not U1784 (N6809,N5758);
not U1785 (N6812,N5762);
buff U1786 (N6815,N5744);
buff U1787 (N6818,N5744);
buff U1788 (N6821,N5755);
buff U1789 (N6824,N5755);
buff U1790 (N6827,N5766);
buff U1791 (N6830,N5766);
and U1792 (N6833,N5850,N5789,N5778,N5771);
and U1793 (N6836,N5771,N3169);
and U1794 (N6837,N5778,N5771,N3173);
and U1795 (N6838,N5789,N5771,N3178,N5778);
and U1796 (N6839,N5778,N3173);
and U1797 (N6840,N5789,N3178,N5778);
and U1798 (N6841,N5850,N5789,N5778);
and U1799 (N6842,N5778,N3173);
and U1800 (N6843,N5789,N3178,N5778);
and U1801 (N6844,N5789,N3178);
and U1802 (N6845,N5856,N5837,N5821,N5807,N5799);
and U1803 (N6848,N5799,N3185);
and U1804 (N6849,N5807,N5799,N3189);
and U1805 (N6850,N5821,N5799,N3195,N5807);
and U1806 (N6851,N5837,N5821,N5799,N3202,N5807);
and U1807 (N6852,N5807,N3189);
and U1808 (N6853,N5821,N3195,N5807);
and U1809 (N6854,N5837,N5821,N3202,N5807);
and U1810 (N6855,N5856,N5821,N5807,N5837);
and U1811 (N6856,N5807,N3189);
and U1812 (N6857,N5821,N3195,N5807);
and U1813 (N6858,N5837,N5821,N3202,N5807);
and U1814 (N6859,N5821,N3195);
and U1815 (N6860,N5837,N5821,N3202);
and U1816 (N6861,N5856,N5821,N5837);
and U1817 (N6862,N5821,N3195);
and U1818 (N6863,N5837,N5821,N3202);
and U1819 (N6864,N5837,N3202);
and U1820 (N6865,N5850,N5789);
and U1821 (N6866,N5856,N5837);
and U1822 (N6867,N5870,N5892,N5881,N5863);
and U1823 (N6870,N5863,N3211);
and U1824 (N6871,N5870,N5863,N3215);
and U1825 (N6872,N5881,N5863,N3221,N5870);
and U1826 (N6873,N5870,N3215);
and U1827 (N6874,N5881,N3221,N5870);
and U1828 (N6875,N5892,N5881,N5870);
and U1829 (N6876,N5870,N3215);
and U1830 (N6877,N3221,N5881,N5870);
and U1831 (N6878,N5881,N3221);
and U1832 (N6879,N5892,N5881);
and U1833 (N6880,N5881,N3221);
and U1834 (N6881,N5905,N5936,N5915,N5898,N5926);
and U1835 (N6884,N5898,N3229);
and U1836 (N6885,N5905,N5898,N3232);
and U1837 (N6886,N5915,N5898,N3236,N5905);
and U1838 (N6887,N5926,N5915,N5898,N3241,N5905);
and U1839 (N6888,N5905,N3232);
and U1840 (N6889,N5915,N3236,N5905);
and U1841 (N6890,N5926,N5915,N3241,N5905);
and U1842 (N6891,N3236,N5915);
and U1843 (N6892,N5926,N5915,N3241);
and U1844 (N6893,N5926,N3241);
nand U1845 (N6894,N5944,N6540);
nand U1846 (N6901,N5946,N6541);
nand U1847 (N6912,N5948,N6542);
nand U1848 (N6923,N5950,N6543);
nand U1849 (N6929,N5952,N6544);
nand U1850 (N6936,N5954,N6545);
nand U1851 (N6946,N5956,N6546);
nand U1852 (N6957,N5958,N6547);
nand U1853 (N6967,N6204,N4575);
not U1854 (N6968,N6204);
not U1855 (N6969,N6207);
nand U1856 (N6970,N5967,N6555);
nand U1857 (N6977,N5969,N6556);
nand U1858 (N6988,N5971,N6557);
nand U1859 (N6998,N5973,N6558);
nand U1860 (N7006,N5975,N6559);
nand U1861 (N7020,N5977,N6560);
nand U1862 (N7036,N5979,N6561);
nand U1863 (N7049,N5989,N6569);
nand U1864 (N7055,N6210,N4610);
not U1865 (N7056,N6210);
and U1866 (N7057,N6021,N6000,N5996,N5991);
and U1867 (N7060,N5991,N3362);
and U1868 (N7061,N5996,N5991,N3363);
and U1869 (N7062,N6000,N5991,N3364,N5996);
and U1870 (N7063,N6022,N6018,N6014,N6009,N6003);
and U1871 (N7064,N6003,N3366);
and U1872 (N7065,N6009,N6003,N3367);
and U1873 (N7066,N6014,N6003,N3368,N6009);
and U1874 (N7067,N6018,N6014,N6003,N3369,N6009);
nand U1875 (N7068,N6594,N6024);
nand U1876 (N7073,N6595,N6026);
nand U1877 (N7077,N6596,N6028);
nand U1878 (N7080,N6597,N6030);
nand U1879 (N7086,N6598,N6599);
nand U1880 (N7091,N6600,N6601);
nand U1881 (N7095,N6602,N6603);
nand U1882 (N7098,N6604,N6038);
nand U1883 (N7099,N6605,N6606);
and U1884 (N7100,N6059,N6056,N6052,N6047,N6041);
and U1885 (N7103,N6041,N3371);
and U1886 (N7104,N6047,N6041,N3372);
and U1887 (N7105,N6052,N6041,N3373,N6047);
and U1888 (N7106,N6056,N6052,N6041,N3374,N6047);
nand U1889 (N7107,N6060,N6621);
nand U1890 (N7114,N6062,N6622);
nand U1891 (N7125,N6064,N6623);
nand U1892 (N7136,N6066,N6624);
nand U1893 (N7142,N6068,N6625);
nand U1894 (N7149,N6070,N6626);
nand U1895 (N7159,N6072,N6627);
nand U1896 (N7170,N6074,N6628);
nand U1897 (N7180,N6076,N6629);
not U1898 (N7187,N6220);
not U1899 (N7188,N6079);
not U1900 (N7191,N6083);
nand U1901 (N7194,N6639,N6091);
nand U1902 (N7198,N6640,N6641);
nand U1903 (N7202,N6642,N6643);
nand U1904 (N7205,N6644,N6097);
nand U1905 (N7209,N6645,N6646);
nand U1906 (N7213,N6647,N6648);
buff U1907 (N7216,N6087);
buff U1908 (N7219,N6087);
nand U1909 (N7222,N6103,N6649);
nand U1910 (N7229,N6105,N6650);
nand U1911 (N7240,N6107,N6651);
nand U1912 (N7250,N6109,N6652);
nand U1913 (N7258,N6111,N6653);
nand U1914 (N7272,N6113,N6654);
nand U1915 (N7288,N6115,N6655);
nand U1916 (N7301,N6117,N6656);
nand U1917 (N7307,N6119,N6657);
nand U1918 (N7314,N6658,N6122);
nand U1919 (N7318,N6659,N6660);
nand U1920 (N7322,N6125,N6661);
not U1921 (N7325,N6127);
not U1922 (N7328,N6131);
nand U1923 (N7331,N6668,N6136);
not U1924 (N7334,N6137);
not U1925 (N7337,N6141);
buff U1926 (N7340,N6145);
buff U1927 (N7343,N6145);
nand U1928 (N7346,N6677,N6678);
nand U1929 (N7351,N6679,N6680);
nand U1930 (N7355,N6681,N6682);
nand U1931 (N7358,N6683,N6684);
nand U1932 (N7364,N6685,N6157);
nand U1933 (N7369,N6686,N6159);
nand U1934 (N7373,N6687,N6161);
nand U1935 (N7376,N6688,N6689);
nand U1936 (N7377,N6164,N6690);
not U1937 (N7378,N6166);
not U1938 (N7381,N6170);
not U1939 (N7384,N6177);
nand U1940 (N7387,N6702,N6703);
nand U1941 (N7391,N6704,N6705);
nand U1942 (N7394,N6706,N6186);
nand U1943 (N7398,N6707,N6708);
nand U1944 (N7402,N6709,N6710);
buff U1945 (N7405,N6174);
buff U1946 (N7408,N6174);
buff U1947 (N7411,N5936);
buff U1948 (N7414,N5898);
buff U1949 (N7417,N5905);
buff U1950 (N7420,N5915);
buff U1951 (N7423,N5926);
buff U1952 (N7426,N5728);
buff U1953 (N7429,N5690);
buff U1954 (N7432,N5697);
buff U1955 (N7435,N5707);
buff U1956 (N7438,N5718);
nand U1957 (N7441,N6192,N6711);
nand U1958 (N7444,N6194,N6712);
buff U1959 (N7447,N5683);
buff U1960 (N7450,N5670);
buff U1961 (N7453,N5632);
buff U1962 (N7456,N5654);
buff U1963 (N7459,N5640);
buff U1964 (N7462,N5640);
buff U1965 (N7465,N5683);
buff U1966 (N7468,N5670);
buff U1967 (N7471,N5632);
buff U1968 (N7474,N5654);
not U1969 (N7477,N6196);
not U1970 (N7478,N6199);
buff U1971 (N7479,N5850);
buff U1972 (N7482,N5789);
buff U1973 (N7485,N5771);
buff U1974 (N7488,N5778);
buff U1975 (N7491,N5850);
buff U1976 (N7494,N5789);
buff U1977 (N7497,N5771);
buff U1978 (N7500,N5778);
buff U1979 (N7503,N5856);
buff U1980 (N7506,N5837);
buff U1981 (N7509,N5799);
buff U1982 (N7512,N5821);
buff U1983 (N7515,N5807);
buff U1984 (N7518,N5807);
buff U1985 (N7521,N5856);
buff U1986 (N7524,N5837);
buff U1987 (N7527,N5799);
buff U1988 (N7530,N5821);
buff U1989 (N7533,N5863);
buff U1990 (N7536,N5863);
buff U1991 (N7539,N5870);
buff U1992 (N7542,N5870);
buff U1993 (N7545,N5881);
buff U1994 (N7548,N5881);
not U1995 (N7551,N6214);
not U1996 (N7552,N6217);
buff U1997 (N7553,N5981);
not U1998 (N7556,N6249);
not U1999 (N7557,N6252);
not U2000 (N7558,N6243);
not U2001 (N7559,N6246);
nand U2002 (N7560,N6731,N6732);
nand U2003 (N7563,N6729,N6730);
nand U2004 (N7566,N6735,N6736);
nand U2005 (N7569,N6733,N6734);
not U2006 (N7572,N6232);
not U2007 (N7573,N6236);
nand U2008 (N7574,N6743,N6744);
nand U2009 (N7577,N6741,N6742);
not U2010 (N7580,N6263);
not U2011 (N7581,N6266);
nand U2012 (N7582,N6753,N6754);
nand U2013 (N7585,N6751,N6752);
nand U2014 (N7588,N6757,N6758);
nand U2015 (N7591,N6755,N6756);
or U2016 (N7609,N3096,N6766,N6767,N6768,N6769);
or U2017 (N7613,N3107,N6782);
or U2018 (N7620,N3136,N6787,N6788,N6789,N6790);
or U2019 (N7649,N3168,N6836,N6837,N6838);
or U2020 (N7650,N3173,N6844);
or U2021 (N7655,N3184,N6848,N6849,N6850,N6851);
or U2022 (N7659,N3195,N6864);
or U2023 (N7668,N3210,N6870,N6871,N6872);
or U2024 (N7671,N3228,N6884,N6885,N6886,N6887);
nand U2025 (N7744,N3661,N6968);
nand U2026 (N7822,N3664,N7056);
or U2027 (N7825,N3361,N7060,N7061,N7062);
or U2028 (N7826,N3365,N7064,N7065,N7066,N7067);
or U2029 (N7852,N3370,N7103,N7104,N7105,N7106);
or U2030 (N8114,N3101,N6777,N6778,N6779);
or U2031 (N8117,N3097,N6770,N6771,N6772,N6773);
nor U2032 (N8131,N3101,N6780,N6781);
nor U2033 (N8134,N3097,N6774,N6775,N6776);
nand U2034 (N8144,N6199,N7477);
nand U2035 (N8145,N6196,N7478);
or U2036 (N8146,N3169,N6839,N6840,N6841);
nor U2037 (N8156,N3169,N6842,N6843);
or U2038 (N8166,N3189,N6859,N6860,N6861);
or U2039 (N8169,N3185,N6852,N6853,N6854,N6855);
nor U2040 (N8183,N3189,N6862,N6863);
nor U2041 (N8186,N3185,N6856,N6857,N6858);
or U2042 (N8196,N3211,N6873,N6874,N6875);
nor U2043 (N8200,N3211,N6876,N6877);
or U2044 (N8204,N3215,N6878,N6879);
nor U2045 (N8208,N3215,N6880);
nand U2046 (N8216,N6252,N7556);
nand U2047 (N8217,N6249,N7557);
nand U2048 (N8218,N6246,N7558);
nand U2049 (N8219,N6243,N7559);
nand U2050 (N8232,N6266,N7580);
nand U2051 (N8233,N6263,N7581);
not U2052 (N8242,N7411);
not U2053 (N8243,N7414);
not U2054 (N8244,N7417);
not U2055 (N8245,N7420);
not U2056 (N8246,N7423);
not U2057 (N8247,N7426);
not U2058 (N8248,N7429);
not U2059 (N8249,N7432);
not U2060 (N8250,N7435);
not U2061 (N8251,N7438);
not U2062 (N8252,N7136);
not U2063 (N8253,N6923);
not U2064 (N8254,N6762);
not U2065 (N8260,N7459);
not U2066 (N8261,N7462);
and U2067 (N8262,N3122,N6762);
and U2068 (N8269,N3155,N6784);
not U2069 (N8274,N6815);
not U2070 (N8275,N6818);
not U2071 (N8276,N6821);
not U2072 (N8277,N6824);
not U2073 (N8278,N6827);
not U2074 (N8279,N6830);
and U2075 (N8280,N5740,N5736,N6815);
and U2076 (N8281,N6800,N6797,N6818);
and U2077 (N8282,N5751,N5747,N6821);
and U2078 (N8283,N6806,N6803,N6824);
and U2079 (N8284,N5762,N5758,N6827);
and U2080 (N8285,N6812,N6809,N6830);
not U2081 (N8288,N6845);
not U2082 (N8294,N7488);
not U2083 (N8295,N7500);
not U2084 (N8296,N7515);
not U2085 (N8297,N7518);
and U2086 (N8298,N6833,N6845);
and U2087 (N8307,N6867,N6881);
not U2088 (N8315,N7533);
not U2089 (N8317,N7536);
not U2090 (N8319,N7539);
not U2091 (N8321,N7542);
nand U2092 (N8322,N7545,N4543);
not U2093 (N8323,N7545);
nand U2094 (N8324,N7548,N5943);
not U2095 (N8325,N7548);
nand U2096 (N8326,N6967,N7744);
and U2097 (N8333,N6901,N6923,N6912,N6894);
and U2098 (N8337,N6894,N4545);
and U2099 (N8338,N6901,N6894,N4549);
and U2100 (N8339,N6912,N6894,N4555,N6901);
and U2101 (N8340,N6901,N4549);
and U2102 (N8341,N6912,N4555,N6901);
and U2103 (N8342,N6923,N6912,N6901);
and U2104 (N8343,N6901,N4549);
and U2105 (N8344,N4555,N6912,N6901);
and U2106 (N8345,N6912,N4555);
and U2107 (N8346,N6923,N6912);
and U2108 (N8347,N6912,N4555);
and U2109 (N8348,N6929,N4563);
and U2110 (N8349,N6936,N6929,N4566);
and U2111 (N8350,N6946,N6929,N4570,N6936);
and U2112 (N8351,N6957,N6946,N6929,N5960,N6936);
and U2113 (N8352,N6936,N4566);
and U2114 (N8353,N6946,N4570,N6936);
and U2115 (N8354,N6957,N6946,N5960,N6936);
and U2116 (N8355,N4570,N6946);
and U2117 (N8356,N6957,N6946,N5960);
and U2118 (N8357,N6957,N5960);
nand U2119 (N8358,N7055,N7822);
and U2120 (N8365,N7049,N6988,N6977,N6970);
and U2121 (N8369,N6970,N4577);
and U2122 (N8370,N6977,N6970,N4581);
and U2123 (N8371,N6988,N6970,N4586,N6977);
and U2124 (N8372,N6977,N4581);
and U2125 (N8373,N6988,N4586,N6977);
and U2126 (N8374,N7049,N6988,N6977);
and U2127 (N8375,N6977,N4581);
and U2128 (N8376,N6988,N4586,N6977);
and U2129 (N8377,N6988,N4586);
and U2130 (N8378,N6998,N4593);
and U2131 (N8379,N7006,N6998,N4597);
and U2132 (N8380,N7020,N6998,N4603,N7006);
and U2133 (N8381,N7036,N7020,N6998,N5981,N7006);
and U2134 (N8382,N7006,N4597);
and U2135 (N8383,N7020,N4603,N7006);
and U2136 (N8384,N7036,N7020,N5981,N7006);
and U2137 (N8385,N7006,N4597);
and U2138 (N8386,N7020,N4603,N7006);
and U2139 (N8387,N7036,N7020,N5981,N7006);
and U2140 (N8388,N7020,N4603);
and U2141 (N8389,N7036,N7020,N5981);
and U2142 (N8390,N7020,N4603);
and U2143 (N8391,N7036,N7020,N5981);
and U2144 (N8392,N7036,N5981);
and U2145 (N8393,N7049,N6988);
and U2146 (N8394,N7057,N7063);
and U2147 (N8404,N7057,N7826);
and U2148 (N8405,N7098,N7077,N7073,N7068);
and U2149 (N8409,N7068,N4632);
and U2150 (N8410,N7073,N7068,N4634);
and U2151 (N8411,N7077,N7068,N4635,N7073);
and U2152 (N8412,N7099,N7095,N7091,N7086,N7080);
and U2153 (N8415,N7080,N4638);
and U2154 (N8416,N7086,N7080,N4639);
and U2155 (N8417,N7091,N7080,N4640,N7086);
and U2156 (N8418,N7095,N7091,N7080,N4641,N7086);
and U2157 (N8421,N3375,N7100);
and U2158 (N8430,N7114,N7136,N7125,N7107);
and U2159 (N8433,N7107,N4657);
and U2160 (N8434,N7114,N7107,N4661);
and U2161 (N8435,N7125,N7107,N4667,N7114);
and U2162 (N8436,N7114,N4661);
and U2163 (N8437,N7125,N4667,N7114);
and U2164 (N8438,N7136,N7125,N7114);
and U2165 (N8439,N7114,N4661);
and U2166 (N8440,N4667,N7125,N7114);
and U2167 (N8441,N7125,N4667);
and U2168 (N8442,N7136,N7125);
and U2169 (N8443,N7125,N4667);
and U2170 (N8444,N7149,N7180,N7159,N7142,N7170);
and U2171 (N8447,N7142,N4675);
and U2172 (N8448,N7149,N7142,N4678);
and U2173 (N8449,N7159,N7142,N4682,N7149);
and U2174 (N8450,N7170,N7159,N7142,N4687,N7149);
and U2175 (N8451,N7149,N4678);
and U2176 (N8452,N7159,N4682,N7149);
and U2177 (N8453,N7170,N7159,N4687,N7149);
and U2178 (N8454,N4682,N7159);
and U2179 (N8455,N7170,N7159,N4687);
and U2180 (N8456,N7170,N4687);
not U2181 (N8457,N7194);
not U2182 (N8460,N7198);
not U2183 (N8463,N7205);
not U2184 (N8466,N7209);
not U2185 (N8469,N7216);
not U2186 (N8470,N7219);
buff U2187 (N8471,N7202);
buff U2188 (N8474,N7202);
buff U2189 (N8477,N7213);
buff U2190 (N8480,N7213);
and U2191 (N8483,N6083,N6079,N7216);
and U2192 (N8484,N7191,N7188,N7219);
and U2193 (N8485,N7301,N7240,N7229,N7222);
and U2194 (N8488,N7222,N4702);
and U2195 (N8489,N7229,N7222,N4706);
and U2196 (N8490,N7240,N7222,N4711,N7229);
and U2197 (N8491,N7229,N4706);
and U2198 (N8492,N7240,N4711,N7229);
and U2199 (N8493,N7301,N7240,N7229);
and U2200 (N8494,N7229,N4706);
and U2201 (N8495,N7240,N4711,N7229);
and U2202 (N8496,N7240,N4711);
and U2203 (N8497,N7307,N7288,N7272,N7258,N7250);
and U2204 (N8500,N7250,N4718);
and U2205 (N8501,N7258,N7250,N4722);
and U2206 (N8502,N7272,N7250,N4728,N7258);
and U2207 (N8503,N7288,N7272,N7250,N4735,N7258);
and U2208 (N8504,N7258,N4722);
and U2209 (N8505,N7272,N4728,N7258);
and U2210 (N8506,N7288,N7272,N4735,N7258);
and U2211 (N8507,N7307,N7272,N7258,N7288);
and U2212 (N8508,N7258,N4722);
and U2213 (N8509,N7272,N4728,N7258);
and U2214 (N8510,N7288,N7272,N4735,N7258);
and U2215 (N8511,N7272,N4728);
and U2216 (N8512,N7288,N7272,N4735);
and U2217 (N8513,N7307,N7272,N7288);
and U2218 (N8514,N7272,N4728);
and U2219 (N8515,N7288,N7272,N4735);
and U2220 (N8516,N7288,N4735);
and U2221 (N8517,N7301,N7240);
and U2222 (N8518,N7307,N7288);
not U2223 (N8519,N7314);
not U2224 (N8522,N7318);
buff U2225 (N8525,N7322);
buff U2226 (N8528,N7322);
buff U2227 (N8531,N7331);
buff U2228 (N8534,N7331);
not U2229 (N8537,N7340);
not U2230 (N8538,N7343);
and U2231 (N8539,N6141,N6137,N7340);
and U2232 (N8540,N7337,N7334,N7343);
and U2233 (N8541,N7376,N7355,N7351,N7346);
and U2234 (N8545,N7346,N4757);
and U2235 (N8546,N7351,N7346,N4758);
and U2236 (N8547,N7355,N7346,N4759,N7351);
and U2237 (N8548,N7377,N7373,N7369,N7364,N7358);
and U2238 (N8551,N7358,N4762);
and U2239 (N8552,N7364,N7358,N4764);
and U2240 (N8553,N7369,N7358,N4766,N7364);
and U2241 (N8554,N7373,N7369,N7358,N4767,N7364);
not U2242 (N8555,N7387);
not U2243 (N8558,N7394);
not U2244 (N8561,N7398);
not U2245 (N8564,N7405);
not U2246 (N8565,N7408);
buff U2247 (N8566,N7391);
buff U2248 (N8569,N7391);
buff U2249 (N8572,N7402);
buff U2250 (N8575,N7402);
and U2251 (N8578,N6170,N6166,N7405);
and U2252 (N8579,N7381,N7378,N7408);
buff U2253 (N8580,N7180);
buff U2254 (N8583,N7142);
buff U2255 (N8586,N7149);
buff U2256 (N8589,N7159);
buff U2257 (N8592,N7170);
buff U2258 (N8595,N6929);
buff U2259 (N8598,N6936);
buff U2260 (N8601,N6946);
buff U2261 (N8604,N6957);
not U2262 (N8607,N7441);
nand U2263 (N8608,N7441,N5469);
not U2264 (N8609,N7444);
nand U2265 (N8610,N7444,N4793);
not U2266 (N8615,N7447);
not U2267 (N8616,N7450);
not U2268 (N8617,N7453);
not U2269 (N8618,N7456);
not U2270 (N8619,N7474);
not U2271 (N8624,N7465);
not U2272 (N8625,N7468);
not U2273 (N8626,N7471);
nand U2274 (N8627,N8144,N8145);
not U2275 (N8632,N7479);
not U2276 (N8633,N7482);
not U2277 (N8634,N7485);
not U2278 (N8637,N7491);
not U2279 (N8638,N7494);
not U2280 (N8639,N7497);
not U2281 (N8644,N7503);
not U2282 (N8645,N7506);
not U2283 (N8646,N7509);
not U2284 (N8647,N7512);
not U2285 (N8648,N7530);
not U2286 (N8653,N7521);
not U2287 (N8654,N7524);
not U2288 (N8655,N7527);
buff U2289 (N8660,N6894);
buff U2290 (N8663,N6894);
buff U2291 (N8666,N6901);
buff U2292 (N8669,N6901);
buff U2293 (N8672,N6912);
buff U2294 (N8675,N6912);
buff U2295 (N8678,N7049);
buff U2296 (N8681,N6988);
buff U2297 (N8684,N6970);
buff U2298 (N8687,N6977);
buff U2299 (N8690,N7049);
buff U2300 (N8693,N6988);
buff U2301 (N8696,N6970);
buff U2302 (N8699,N6977);
buff U2303 (N8702,N7036);
buff U2304 (N8705,N6998);
buff U2305 (N8708,N7020);
buff U2306 (N8711,N7006);
buff U2307 (N8714,N7006);
not U2308 (N8717,N7553);
buff U2309 (N8718,N7036);
buff U2310 (N8721,N6998);
buff U2311 (N8724,N7020);
nand U2312 (N8727,N8216,N8217);
nand U2313 (N8730,N8218,N8219);
not U2314 (N8733,N7574);
not U2315 (N8734,N7577);
buff U2316 (N8735,N7107);
buff U2317 (N8738,N7107);
buff U2318 (N8741,N7114);
buff U2319 (N8744,N7114);
buff U2320 (N8747,N7125);
buff U2321 (N8750,N7125);
not U2322 (N8753,N7560);
not U2323 (N8754,N7563);
not U2324 (N8755,N7566);
not U2325 (N8756,N7569);
buff U2326 (N8757,N7301);
buff U2327 (N8760,N7240);
buff U2328 (N8763,N7222);
buff U2329 (N8766,N7229);
buff U2330 (N8769,N7301);
buff U2331 (N8772,N7240);
buff U2332 (N8775,N7222);
buff U2333 (N8778,N7229);
buff U2334 (N8781,N7307);
buff U2335 (N8784,N7288);
buff U2336 (N8787,N7250);
buff U2337 (N8790,N7272);
buff U2338 (N8793,N7258);
buff U2339 (N8796,N7258);
buff U2340 (N8799,N7307);
buff U2341 (N8802,N7288);
buff U2342 (N8805,N7250);
buff U2343 (N8808,N7272);
nand U2344 (N8811,N8232,N8233);
not U2345 (N8814,N7588);
not U2346 (N8815,N7591);
not U2347 (N8816,N7582);
not U2348 (N8817,N7585);
and U2349 (N8818,N7620,N3155);
and U2350 (N8840,N3122,N7609);
not U2351 (N8857,N7609);
and U2352 (N8861,N6797,N5740,N8274);
and U2353 (N8862,N5736,N6800,N8275);
and U2354 (N8863,N6803,N5751,N8276);
and U2355 (N8864,N5747,N6806,N8277);
and U2356 (N8865,N6809,N5762,N8278);
and U2357 (N8866,N5758,N6812,N8279);
not U2358 (N8871,N7655);
and U2359 (N8874,N6833,N7655);
and U2360 (N8878,N7671,N6867);
not U2361 (N8879,N8196);
nand U2362 (N8880,N8196,N8315);
not U2363 (N8881,N8200);
nand U2364 (N8882,N8200,N8317);
not U2365 (N8883,N8204);
nand U2366 (N8884,N8204,N8319);
not U2367 (N8885,N8208);
nand U2368 (N8886,N8208,N8321);
nand U2369 (N8887,N3658,N8323);
nand U2370 (N8888,N4817,N8325);
or U2371 (N8898,N4544,N8337,N8338,N8339);
or U2372 (N8902,N4562,N8348,N8349,N8350,N8351);
or U2373 (N8920,N4576,N8369,N8370,N8371);
or U2374 (N8924,N4581,N8377);
or U2375 (N8927,N4592,N8378,N8379,N8380,N8381);
or U2376 (N8931,N4603,N8392);
or U2377 (N8943,N7825,N8404);
or U2378 (N8950,N4630,N8409,N8410,N8411);
or U2379 (N8956,N4637,N8415,N8416,N8417,N8418);
not U2380 (N8959,N7852);
and U2381 (N8960,N3375,N7852);
or U2382 (N8963,N4656,N8433,N8434,N8435);
or U2383 (N8966,N4674,N8447,N8448,N8449,N8450);
and U2384 (N8991,N7188,N6083,N8469);
and U2385 (N8992,N6079,N7191,N8470);
or U2386 (N8995,N4701,N8488,N8489,N8490);
or U2387 (N8996,N4706,N8496);
or U2388 (N9001,N4717,N8500,N8501,N8502,N8503);
or U2389 (N9005,N4728,N8516);
and U2390 (N9024,N7334,N6141,N8537);
and U2391 (N9025,N6137,N7337,N8538);
or U2392 (N9029,N4756,N8545,N8546,N8547);
or U2393 (N9035,N4760,N8551,N8552,N8553,N8554);
and U2394 (N9053,N7378,N6170,N8564);
and U2395 (N9054,N6166,N7381,N8565);
nand U2396 (N9064,N4303,N8607);
nand U2397 (N9065,N3507,N8609);
not U2398 (N9066,N8114);
nand U2399 (N9067,N8114,N4795);
or U2400 (N9068,N7613,N6783);
not U2401 (N9071,N8117);
not U2402 (N9072,N8131);
nand U2403 (N9073,N8131,N6195);
not U2404 (N9074,N7613);
not U2405 (N9077,N8134);
or U2406 (N9079,N7650,N6865);
not U2407 (N9082,N8146);
not U2408 (N9083,N7650);
not U2409 (N9086,N8156);
not U2410 (N9087,N8166);
nand U2411 (N9088,N8166,N4813);
or U2412 (N9089,N7659,N6866);
not U2413 (N9092,N8169);
not U2414 (N9093,N8183);
nand U2415 (N9094,N8183,N6203);
not U2416 (N9095,N7659);
not U2417 (N9098,N8186);
or U2418 (N9099,N4545,N8340,N8341,N8342);
nor U2419 (N9103,N4545,N8343,N8344);
or U2420 (N9107,N4549,N8345,N8346);
nor U2421 (N9111,N4549,N8347);
or U2422 (N9117,N4577,N8372,N8373,N8374);
nor U2423 (N9127,N4577,N8375,N8376);
nor U2424 (N9146,N4597,N8390,N8391);
nor U2425 (N9149,N4593,N8385,N8386,N8387);
nand U2426 (N9159,N7577,N8733);
nand U2427 (N9160,N7574,N8734);
or U2428 (N9161,N4657,N8436,N8437,N8438);
nor U2429 (N9165,N4657,N8439,N8440);
or U2430 (N9169,N4661,N8441,N8442);
nor U2431 (N9173,N4661,N8443);
nand U2432 (N9179,N7563,N8753);
nand U2433 (N9180,N7560,N8754);
nand U2434 (N9181,N7569,N8755);
nand U2435 (N9182,N7566,N8756);
or U2436 (N9183,N4702,N8491,N8492,N8493);
nor U2437 (N9193,N4702,N8494,N8495);
or U2438 (N9203,N4722,N8511,N8512,N8513);
or U2439 (N9206,N4718,N8504,N8505,N8506,N8507);
nor U2440 (N9220,N4722,N8514,N8515);
nor U2441 (N9223,N4718,N8508,N8509,N8510);
nand U2442 (N9234,N7591,N8814);
nand U2443 (N9235,N7588,N8815);
nand U2444 (N9236,N7585,N8816);
nand U2445 (N9237,N7582,N8817);
or U2446 (N9238,N3159,N8818);
or U2447 (N9242,N3126,N8840);
nand U2448 (N9243,N8324,N8888);
not U2449 (N9244,N8580);
not U2450 (N9245,N8583);
not U2451 (N9246,N8586);
not U2452 (N9247,N8589);
not U2453 (N9248,N8592);
not U2454 (N9249,N8595);
not U2455 (N9250,N8598);
not U2456 (N9251,N8601);
not U2457 (N9252,N8604);
nor U2458 (N9256,N8861,N8280);
nor U2459 (N9257,N8862,N8281);
nor U2460 (N9258,N8863,N8282);
nor U2461 (N9259,N8864,N8283);
nor U2462 (N9260,N8865,N8284);
nor U2463 (N9261,N8866,N8285);
not U2464 (N9262,N8627);
or U2465 (N9265,N7649,N8874);
or U2466 (N9268,N7668,N8878);
nand U2467 (N9271,N7533,N8879);
nand U2468 (N9272,N7536,N8881);
nand U2469 (N9273,N7539,N8883);
nand U2470 (N9274,N7542,N8885);
nand U2471 (N9275,N8322,N8887);
not U2472 (N9276,N8333);
and U2473 (N9280,N6936,N8326,N6946,N6929,N6957);
and U2474 (N9285,N367,N8326,N6946,N6957,N6936);
and U2475 (N9286,N367,N8326,N6946,N6957);
and U2476 (N9287,N367,N8326,N6957);
and U2477 (N9288,N367,N8326);
not U2478 (N9290,N8660);
not U2479 (N9292,N8663);
not U2480 (N9294,N8666);
not U2481 (N9296,N8669);
nand U2482 (N9297,N8672,N5966);
not U2483 (N9298,N8672);
nand U2484 (N9299,N8675,N6969);
not U2485 (N9300,N8675);
not U2486 (N9301,N8365);
and U2487 (N9307,N8358,N7036,N7020,N7006,N6998);
and U2488 (N9314,N8358,N7020,N7006,N7036);
and U2489 (N9315,N8358,N7020,N7036);
and U2490 (N9318,N8358,N7036);
not U2491 (N9319,N8687);
not U2492 (N9320,N8699);
not U2493 (N9321,N8711);
not U2494 (N9322,N8714);
not U2495 (N9323,N8727);
not U2496 (N9324,N8730);
not U2497 (N9326,N8405);
and U2498 (N9332,N8405,N8412);
or U2499 (N9339,N4193,N8960);
and U2500 (N9344,N8430,N8444);
not U2501 (N9352,N8735);
not U2502 (N9354,N8738);
not U2503 (N9356,N8741);
not U2504 (N9358,N8744);
nand U2505 (N9359,N8747,N6078);
not U2506 (N9360,N8747);
nand U2507 (N9361,N8750,N7187);
not U2508 (N9362,N8750);
not U2509 (N9363,N8471);
not U2510 (N9364,N8474);
not U2511 (N9365,N8477);
not U2512 (N9366,N8480);
nor U2513 (N9367,N8991,N8483);
nor U2514 (N9368,N8992,N8484);
and U2515 (N9369,N7198,N7194,N8471);
and U2516 (N9370,N8460,N8457,N8474);
and U2517 (N9371,N7209,N7205,N8477);
and U2518 (N9372,N8466,N8463,N8480);
not U2519 (N9375,N8497);
not U2520 (N9381,N8766);
not U2521 (N9382,N8778);
not U2522 (N9383,N8793);
not U2523 (N9384,N8796);
and U2524 (N9385,N8485,N8497);
not U2525 (N9392,N8525);
not U2526 (N9393,N8528);
not U2527 (N9394,N8531);
not U2528 (N9395,N8534);
and U2529 (N9396,N7318,N7314,N8525);
and U2530 (N9397,N8522,N8519,N8528);
and U2531 (N9398,N6131,N6127,N8531);
and U2532 (N9399,N7328,N7325,N8534);
nor U2533 (N9400,N9024,N8539);
nor U2534 (N9401,N9025,N8540);
not U2535 (N9402,N8541);
nand U2536 (N9407,N8548,N89);
and U2537 (N9408,N8541,N8548);
not U2538 (N9412,N8811);
not U2539 (N9413,N8566);
not U2540 (N9414,N8569);
not U2541 (N9415,N8572);
not U2542 (N9416,N8575);
nor U2543 (N9417,N9053,N8578);
nor U2544 (N9418,N9054,N8579);
and U2545 (N9419,N7387,N6177,N8566);
and U2546 (N9420,N8555,N7384,N8569);
and U2547 (N9421,N7398,N7394,N8572);
and U2548 (N9422,N8561,N8558,N8575);
buff U2549 (N9423,N8326);
nand U2550 (N9426,N9064,N8608);
nand U2551 (N9429,N9065,N8610);
nand U2552 (N9432,N3515,N9066);
nand U2553 (N9435,N4796,N9072);
nand U2554 (N9442,N3628,N9087);
nand U2555 (N9445,N4814,N9093);
not U2556 (N9454,N8678);
not U2557 (N9455,N8681);
not U2558 (N9456,N8684);
not U2559 (N9459,N8690);
not U2560 (N9460,N8693);
not U2561 (N9461,N8696);
buff U2562 (N9462,N8358);
not U2563 (N9465,N8702);
not U2564 (N9466,N8705);
not U2565 (N9467,N8708);
not U2566 (N9468,N8724);
buff U2567 (N9473,N8358);
not U2568 (N9476,N8718);
not U2569 (N9477,N8721);
nand U2570 (N9478,N9159,N9160);
nand U2571 (N9485,N9179,N9180);
nand U2572 (N9488,N9181,N9182);
not U2573 (N9493,N8757);
not U2574 (N9494,N8760);
not U2575 (N9495,N8763);
not U2576 (N9498,N8769);
not U2577 (N9499,N8772);
not U2578 (N9500,N8775);
not U2579 (N9505,N8781);
not U2580 (N9506,N8784);
not U2581 (N9507,N8787);
not U2582 (N9508,N8790);
not U2583 (N9509,N8808);
not U2584 (N9514,N8799);
not U2585 (N9515,N8802);
not U2586 (N9516,N8805);
nand U2587 (N9517,N9234,N9235);
nand U2588 (N9520,N9236,N9237);
and U2589 (N9526,N8943,N8421);
and U2590 (N9531,N8943,N8421);
nand U2591 (N9539,N9271,N8880);
nand U2592 (N9540,N9273,N8884);
not U2593 (N9541,N9275);
and U2594 (N9543,N8857,N8254);
and U2595 (N9551,N8871,N8288);
nand U2596 (N9555,N9272,N8882);
nand U2597 (N9556,N9274,N8886);
not U2598 (N9557,N8898);
and U2599 (N9560,N8902,N8333);
not U2600 (N9561,N9099);
nand U2601 (N9562,N9099,N9290);
not U2602 (N9563,N9103);
nand U2603 (N9564,N9103,N9292);
not U2604 (N9565,N9107);
nand U2605 (N9566,N9107,N9294);
not U2606 (N9567,N9111);
nand U2607 (N9568,N9111,N9296);
nand U2608 (N9569,N4844,N9298);
nand U2609 (N9570,N6207,N9300);
not U2610 (N9571,N8920);
not U2611 (N9575,N8927);
and U2612 (N9579,N8365,N8927);
not U2613 (N9581,N8950);
not U2614 (N9582,N8956);
and U2615 (N9585,N8405,N8956);
and U2616 (N9591,N8966,N8430);
not U2617 (N9592,N9161);
nand U2618 (N9593,N9161,N9352);
not U2619 (N9594,N9165);
nand U2620 (N9595,N9165,N9354);
not U2621 (N9596,N9169);
nand U2622 (N9597,N9169,N9356);
not U2623 (N9598,N9173);
nand U2624 (N9599,N9173,N9358);
nand U2625 (N9600,N4940,N9360);
nand U2626 (N9601,N6220,N9362);
and U2627 (N9602,N8457,N7198,N9363);
and U2628 (N9603,N7194,N8460,N9364);
and U2629 (N9604,N8463,N7209,N9365);
and U2630 (N9605,N7205,N8466,N9366);
not U2631 (N9608,N9001);
and U2632 (N9611,N8485,N9001);
and U2633 (N9612,N8519,N7318,N9392);
and U2634 (N9613,N7314,N8522,N9393);
and U2635 (N9614,N7325,N6131,N9394);
and U2636 (N9615,N6127,N7328,N9395);
not U2637 (N9616,N9029);
not U2638 (N9617,N9035);
and U2639 (N9618,N8541,N9035);
and U2640 (N9621,N7384,N7387,N9413);
and U2641 (N9622,N6177,N8555,N9414);
and U2642 (N9623,N8558,N7398,N9415);
and U2643 (N9624,N7394,N8561,N9416);
or U2644 (N9626,N4563,N8352,N8353,N8354,N9285);
or U2645 (N9629,N4566,N8355,N8356,N9286);
or U2646 (N9632,N4570,N8357,N9287);
or U2647 (N9635,N5960,N9288);
nand U2648 (N9642,N9067,N9432);
not U2649 (N9645,N9068);
nand U2650 (N9646,N9073,N9435);
not U2651 (N9649,N9074);
nand U2652 (N9650,N9257,N9256);
nand U2653 (N9653,N9259,N9258);
nand U2654 (N9656,N9261,N9260);
not U2655 (N9659,N9079);
nand U2656 (N9660,N9079,N4809);
not U2657 (N9661,N9083);
nand U2658 (N9662,N9083,N6202);
nand U2659 (N9663,N9088,N9442);
not U2660 (N9666,N9089);
nand U2661 (N9667,N9094,N9445);
not U2662 (N9670,N9095);
or U2663 (N9671,N8924,N8393);
not U2664 (N9674,N9117);
not U2665 (N9675,N8924);
not U2666 (N9678,N9127);
or U2667 (N9679,N4597,N8388,N8389,N9315);
or U2668 (N9682,N8931,N9318);
or U2669 (N9685,N4593,N8382,N8383,N8384,N9314);
not U2670 (N9690,N9146);
nand U2671 (N9691,N9146,N8717);
not U2672 (N9692,N8931);
not U2673 (N9695,N9149);
nand U2674 (N9698,N9401,N9400);
nand U2675 (N9702,N9368,N9367);
or U2676 (N9707,N8996,N8517);
not U2677 (N9710,N9183);
not U2678 (N9711,N8996);
not U2679 (N9714,N9193);
not U2680 (N9715,N9203);
nand U2681 (N9716,N9203,N6235);
or U2682 (N9717,N9005,N8518);
not U2683 (N9720,N9206);
not U2684 (N9721,N9220);
nand U2685 (N9722,N9220,N7573);
not U2686 (N9723,N9005);
not U2687 (N9726,N9223);
nand U2688 (N9727,N9418,N9417);
and U2689 (N9732,N9268,N8269);
nand U2690 (N9733,N9581,N9326);
and U2691 (N9734,N89,N9408,N9332,N8394,N8421);
and U2692 (N9735,N89,N9408,N9332,N8394,N8421);
and U2693 (N9736,N9265,N8262);
not U2694 (N9737,N9555);
not U2695 (N9738,N9556);
nand U2696 (N9739,N9361,N9601);
nand U2697 (N9740,N9423,N1115);
not U2698 (N9741,N9423);
nand U2699 (N9742,N9299,N9570);
and U2700 (N9754,N8333,N9280);
or U2701 (N9758,N8898,N9560);
nand U2702 (N9762,N8660,N9561);
nand U2703 (N9763,N8663,N9563);
nand U2704 (N9764,N8666,N9565);
nand U2705 (N9765,N8669,N9567);
nand U2706 (N9766,N9297,N9569);
and U2707 (N9767,N9280,N367);
nand U2708 (N9768,N9557,N9276);
not U2709 (N9769,N9307);
nand U2710 (N9773,N9307,N367);
nand U2711 (N9774,N9571,N9301);
and U2712 (N9775,N8365,N9307);
or U2713 (N9779,N8920,N9579);
not U2714 (N9784,N9478);
nand U2715 (N9785,N9616,N9402);
or U2716 (N9786,N8950,N9585);
and U2717 (N9790,N89,N9408,N9332,N8394);
or U2718 (N9791,N8963,N9591);
nand U2719 (N9795,N8735,N9592);
nand U2720 (N9796,N8738,N9594);
nand U2721 (N9797,N8741,N9596);
nand U2722 (N9798,N8744,N9598);
nand U2723 (N9799,N9359,N9600);
nor U2724 (N9800,N9602,N9369);
nor U2725 (N9801,N9603,N9370);
nor U2726 (N9802,N9604,N9371);
nor U2727 (N9803,N9605,N9372);
not U2728 (N9805,N9485);
not U2729 (N9806,N9488);
or U2730 (N9809,N8995,N9611);
nor U2731 (N9813,N9612,N9396);
nor U2732 (N9814,N9613,N9397);
nor U2733 (N9815,N9614,N9398);
nor U2734 (N9816,N9615,N9399);
and U2735 (N9817,N9617,N9407);
or U2736 (N9820,N9029,N9618);
not U2737 (N9825,N9517);
not U2738 (N9826,N9520);
nor U2739 (N9827,N9621,N9419);
nor U2740 (N9828,N9622,N9420);
nor U2741 (N9829,N9623,N9421);
nor U2742 (N9830,N9624,N9422);
not U2743 (N9835,N9426);
nand U2744 (N9836,N9426,N4789);
not U2745 (N9837,N9429);
nand U2746 (N9838,N9429,N4794);
nand U2747 (N9846,N3625,N9659);
nand U2748 (N9847,N4810,N9661);
not U2749 (N9862,N9462);
nand U2750 (N9863,N7553,N9690);
not U2751 (N9866,N9473);
nand U2752 (N9873,N5030,N9715);
nand U2753 (N9876,N6236,N9721);
nand U2754 (N9890,N9795,N9593);
nand U2755 (N9891,N9797,N9597);
not U2756 (N9892,N9799);
nand U2757 (N9893,N871,N9741);
nand U2758 (N9894,N9762,N9562);
nand U2759 (N9895,N9764,N9566);
not U2760 (N9896,N9766);
not U2761 (N9897,N9626);
nand U2762 (N9898,N9626,N9249);
not U2763 (N9899,N9629);
nand U2764 (N9900,N9629,N9250);
not U2765 (N9901,N9632);
nand U2766 (N9902,N9632,N9251);
not U2767 (N9903,N9635);
nand U2768 (N9904,N9635,N9252);
not U2769 (N9905,N9543);
not U2770 (N9906,N9650);
nand U2771 (N9907,N9650,N5769);
not U2772 (N9908,N9653);
nand U2773 (N9909,N9653,N5770);
not U2774 (N9910,N9656);
nand U2775 (N9911,N9656,N9262);
not U2776 (N9917,N9551);
nand U2777 (N9923,N9763,N9564);
nand U2778 (N9924,N9765,N9568);
or U2779 (N9925,N8902,N9767);
and U2780 (N9932,N9575,N9773);
and U2781 (N9935,N9575,N9769);
not U2782 (N9938,N9698);
nand U2783 (N9939,N9698,N9323);
nand U2784 (N9945,N9796,N9595);
nand U2785 (N9946,N9798,N9599);
not U2786 (N9947,N9702);
nand U2787 (N9948,N9702,N6102);
and U2788 (N9949,N9608,N9375);
not U2789 (N9953,N9727);
nand U2790 (N9954,N9727,N9412);
nand U2791 (N9955,N3502,N9835);
nand U2792 (N9956,N3510,N9837);
not U2793 (N9957,N9642);
nand U2794 (N9958,N9642,N9645);
not U2795 (N9959,N9646);
nand U2796 (N9960,N9646,N9649);
nand U2797 (N9961,N9660,N9846);
nand U2798 (N9964,N9662,N9847);
not U2799 (N9967,N9663);
nand U2800 (N9968,N9663,N9666);
not U2801 (N9969,N9667);
nand U2802 (N9970,N9667,N9670);
not U2803 (N9971,N9671);
nand U2804 (N9972,N9671,N6213);
not U2805 (N9973,N9675);
nand U2806 (N9974,N9675,N7551);
not U2807 (N9975,N9679);
nand U2808 (N9976,N9679,N7552);
not U2809 (N9977,N9682);
not U2810 (N9978,N9685);
nand U2811 (N9979,N9691,N9863);
not U2812 (N9982,N9692);
nand U2813 (N9983,N9814,N9813);
nand U2814 (N9986,N9816,N9815);
nand U2815 (N9989,N9801,N9800);
nand U2816 (N9992,N9803,N9802);
not U2817 (N9995,N9707);
nand U2818 (N9996,N9707,N6231);
not U2819 (N9997,N9711);
nand U2820 (N9998,N9711,N7572);
nand U2821 (N9999,N9716,N9873);
not U2822 (N10002,N9717);
nand U2823 (N10003,N9722,N9876);
not U2824 (N10006,N9723);
nand U2825 (N10007,N9830,N9829);
nand U2826 (N10010,N9828,N9827);
and U2827 (N10013,N9791,N8307,N8269);
and U2828 (N10014,N9758,N9344,N8307,N8269);
and U2829 (N10015,N367,N9754,N9344,N8307,N8269);
and U2830 (N10016,N9786,N8394,N8421);
and U2831 (N10017,N9820,N9332,N8394,N8421);
and U2832 (N10018,N9786,N8394,N8421);
and U2833 (N10019,N9820,N9332,N8394,N8421);
and U2834 (N10020,N9809,N8298,N8262);
and U2835 (N10021,N9779,N9385,N8298,N8262);
and U2836 (N10022,N367,N9775,N9385,N8298,N8262);
not U2837 (N10023,N9945);
not U2838 (N10024,N9946);
nand U2839 (N10025,N9740,N9893);
not U2840 (N10026,N9923);
not U2841 (N10028,N9924);
nand U2842 (N10032,N8595,N9897);
nand U2843 (N10033,N8598,N9899);
nand U2844 (N10034,N8601,N9901);
nand U2845 (N10035,N8604,N9903);
nand U2846 (N10036,N4803,N9906);
nand U2847 (N10037,N4806,N9908);
nand U2848 (N10038,N8627,N9910);
and U2849 (N10039,N9809,N8298);
and U2850 (N10040,N9779,N9385,N8298);
and U2851 (N10041,N367,N9775,N9385,N8298);
and U2852 (N10042,N9779,N9385);
and U2853 (N10043,N367,N9775,N9385);
nand U2854 (N10050,N8727,N9938);
not U2855 (N10053,N9817);
and U2856 (N10054,N9817,N9029);
and U2857 (N10055,N9786,N8394);
and U2858 (N10056,N9820,N9332,N8394);
and U2859 (N10057,N9791,N8307);
and U2860 (N10058,N9758,N9344,N8307);
and U2861 (N10059,N367,N9754,N9344,N8307);
and U2862 (N10060,N9758,N9344);
and U2863 (N10061,N367,N9754,N9344);
nand U2864 (N10062,N4997,N9947);
nand U2865 (N10067,N8811,N9953);
nand U2866 (N10070,N9955,N9836);
nand U2867 (N10073,N9956,N9838);
nand U2868 (N10076,N9068,N9957);
nand U2869 (N10077,N9074,N9959);
nand U2870 (N10082,N9089,N9967);
nand U2871 (N10083,N9095,N9969);
nand U2872 (N10084,N4871,N9971);
nand U2873 (N10085,N6214,N9973);
nand U2874 (N10086,N6217,N9975);
nand U2875 (N10093,N5027,N9995);
nand U2876 (N10094,N6232,N9997);
or U2877 (N10101,N9238,N9732,N10013,N10014,N10015);
or U2878 (N10102,N9339,N9526,N10016,N10017,N9734);
or U2879 (N10103,N9339,N9531,N10018,N10019,N9735);
or U2880 (N10104,N9242,N9736,N10020,N10021,N10022);
and U2881 (N10105,N9925,N9894);
and U2882 (N10106,N9925,N9895);
and U2883 (N10107,N9925,N9896);
and U2884 (N10108,N9925,N8253);
nand U2885 (N10109,N10032,N9898);
nand U2886 (N10110,N10033,N9900);
nand U2887 (N10111,N10034,N9902);
nand U2888 (N10112,N10035,N9904);
nand U2889 (N10113,N10036,N9907);
nand U2890 (N10114,N10037,N9909);
nand U2891 (N10115,N10038,N9911);
or U2892 (N10116,N9265,N10039,N10040,N10041);
or U2893 (N10119,N9809,N10042,N10043);
not U2894 (N10124,N9925);
and U2895 (N10130,N9768,N9925);
not U2896 (N10131,N9932);
not U2897 (N10132,N9935);
and U2898 (N10133,N9932,N8920);
nand U2899 (N10134,N10050,N9939);
not U2900 (N10135,N9983);
nand U2901 (N10136,N9983,N9324);
not U2902 (N10137,N9986);
nand U2903 (N10138,N9986,N9784);
and U2904 (N10139,N9785,N10053);
or U2905 (N10140,N8943,N10055,N10056,N9790);
or U2906 (N10141,N9268,N10057,N10058,N10059);
or U2907 (N10148,N9791,N10060,N10061);
nand U2908 (N10155,N10062,N9948);
not U2909 (N10156,N9989);
nand U2910 (N10157,N9989,N9805);
not U2911 (N10158,N9992);
nand U2912 (N10159,N9992,N9806);
not U2913 (N10160,N9949);
nand U2914 (N10161,N10067,N9954);
not U2915 (N10162,N10007);
nand U2916 (N10163,N10007,N9825);
not U2917 (N10164,N10010);
nand U2918 (N10165,N10010,N9826);
nand U2919 (N10170,N10076,N9958);
nand U2920 (N10173,N10077,N9960);
not U2921 (N10176,N9961);
nand U2922 (N10177,N9961,N9082);
not U2923 (N10178,N9964);
nand U2924 (N10179,N9964,N9086);
nand U2925 (N10180,N10082,N9968);
nand U2926 (N10183,N10083,N9970);
nand U2927 (N10186,N9972,N10084);
nand U2928 (N10189,N9974,N10085);
nand U2929 (N10192,N9976,N10086);
not U2930 (N10195,N9979);
nand U2931 (N10196,N9979,N9982);
nand U2932 (N10197,N9996,N10093);
nand U2933 (N10200,N9998,N10094);
not U2934 (N10203,N9999);
nand U2935 (N10204,N9999,N10002);
not U2936 (N10205,N10003);
nand U2937 (N10206,N10003,N10006);
nand U2938 (N10212,N10070,N4308);
nand U2939 (N10213,N10073,N4313);
and U2940 (N10230,N9774,N10131);
nand U2941 (N10231,N8730,N10135);
nand U2942 (N10232,N9478,N10137);
or U2943 (N10233,N10139,N10054);
nand U2944 (N10234,N7100,N10140);
nand U2945 (N10237,N9485,N10156);
nand U2946 (N10238,N9488,N10158);
nand U2947 (N10239,N9517,N10162);
nand U2948 (N10240,N9520,N10164);
not U2949 (N10241,N10070);
not U2950 (N10242,N10073);
nand U2951 (N10247,N8146,N10176);
nand U2952 (N10248,N8156,N10178);
nand U2953 (N10259,N9692,N10195);
nand U2954 (N10264,N9717,N10203);
nand U2955 (N10265,N9723,N10205);
and U2956 (N10266,N10026,N10124);
and U2957 (N10267,N10028,N10124);
and U2958 (N10268,N9742,N10124);
and U2959 (N10269,N6923,N10124);
nand U2960 (N10270,N6762,N10116);
nand U2961 (N10271,N3061,N10241);
nand U2962 (N10272,N3064,N10242);
buff U2963 (N10273,N10116);
and U2964 (N10278,N10141,N5728,N5707,N5718,N5697);
and U2965 (N10279,N10141,N5728,N5707,N5718);
and U2966 (N10280,N10141,N5728,N5718);
and U2967 (N10281,N10141,N5728);
and U2968 (N10282,N6784,N10141);
not U2969 (N10283,N10119);
and U2970 (N10287,N10148,N5936,N5915,N5926,N5905);
and U2971 (N10288,N10148,N5936,N5915,N5926);
and U2972 (N10289,N10148,N5936,N5926);
and U2973 (N10290,N10148,N5936);
and U2974 (N10291,N6881,N10148);
and U2975 (N10292,N8898,N10124);
nand U2976 (N10293,N10231,N10136);
nand U2977 (N10294,N10232,N10138);
nand U2978 (N10295,N8412,N10233);
and U2979 (N10296,N8959,N10234);
nand U2980 (N10299,N10237,N10157);
nand U2981 (N10300,N10238,N10159);
or U2982 (N10301,N10230,N10133);
nand U2983 (N10306,N10239,N10163);
nand U2984 (N10307,N10240,N10165);
buff U2985 (N10308,N10148);
buff U2986 (N10311,N10141);
not U2987 (N10314,N10170);
nand U2988 (N10315,N10170,N9071);
not U2989 (N10316,N10173);
nand U2990 (N10317,N10173,N9077);
nand U2991 (N10318,N10247,N10177);
nand U2992 (N10321,N10248,N10179);
not U2993 (N10324,N10180);
nand U2994 (N10325,N10180,N9092);
not U2995 (N10326,N10183);
nand U2996 (N10327,N10183,N9098);
not U2997 (N10328,N10186);
nand U2998 (N10329,N10186,N9674);
not U2999 (N10330,N10189);
nand U3000 (N10331,N10189,N9678);
not U3001 (N10332,N10192);
nand U3002 (N10333,N10192,N9977);
nand U3003 (N10334,N10259,N10196);
not U3004 (N10337,N10197);
nand U3005 (N10338,N10197,N9710);
not U3006 (N10339,N10200);
nand U3007 (N10340,N10200,N9714);
nand U3008 (N10341,N10264,N10204);
nand U3009 (N10344,N10265,N10206);
or U3010 (N10350,N10266,N10105);
or U3011 (N10351,N10267,N10106);
or U3012 (N10352,N10268,N10107);
or U3013 (N10353,N10269,N10108);
and U3014 (N10354,N8857,N10270);
nand U3015 (N10357,N10271,N10212);
nand U3016 (N10360,N10272,N10213);
or U3017 (N10367,N7620,N10282);
or U3018 (N10375,N7671,N10291);
or U3019 (N10381,N10292,N10130);
and U3020 (N10388,N10114,N10134,N10293,N10294);
and U3021 (N10391,N9582,N10295);
and U3022 (N10399,N10113,N10115,N10299,N10300);
and U3023 (N10402,N10155,N10161,N10306,N10307);
or U3024 (N10406,N3229,N6888,N6889,N6890,N10287);
or U3025 (N10409,N3232,N6891,N6892,N10288);
or U3026 (N10412,N3236,N6893,N10289);
or U3027 (N10415,N3241,N10290);
or U3028 (N10419,N3137,N6791,N6792,N6793,N10278);
or U3029 (N10422,N3140,N6794,N6795,N10279);
or U3030 (N10425,N3144,N6796,N10280);
or U3031 (N10428,N3149,N10281);
nand U3032 (N10431,N8117,N10314);
nand U3033 (N10432,N8134,N10316);
nand U3034 (N10437,N8169,N10324);
nand U3035 (N10438,N8186,N10326);
nand U3036 (N10439,N9117,N10328);
nand U3037 (N10440,N9127,N10330);
nand U3038 (N10441,N9682,N10332);
nand U3039 (N10444,N9183,N10337);
nand U3040 (N10445,N9193,N10339);
not U3041 (N10450,N10296);
and U3042 (N10451,N10296,N4193);
not U3043 (N10455,N10308);
nand U3044 (N10456,N10308,N8242);
not U3045 (N10465,N10311);
nand U3046 (N10466,N10311,N8247);
not U3047 (N10479,N10273);
not U3048 (N10497,N10301);
nand U3049 (N10509,N10431,N10315);
nand U3050 (N10512,N10432,N10317);
not U3051 (N10515,N10318);
nand U3052 (N10516,N10318,N8632);
not U3053 (N10517,N10321);
nand U3054 (N10518,N10321,N8637);
nand U3055 (N10519,N10437,N10325);
nand U3056 (N10522,N10438,N10327);
nand U3057 (N10525,N10439,N10329);
nand U3058 (N10528,N10440,N10331);
nand U3059 (N10531,N10441,N10333);
not U3060 (N10534,N10334);
nand U3061 (N10535,N10334,N9695);
nand U3062 (N10536,N10444,N10338);
nand U3063 (N10539,N10445,N10340);
not U3064 (N10542,N10341);
nand U3065 (N10543,N10341,N9720);
not U3066 (N10544,N10344);
nand U3067 (N10545,N10344,N9726);
and U3068 (N10546,N5631,N10450);
not U3069 (N10547,N10391);
and U3070 (N10548,N10391,N8950);
and U3071 (N10549,N5165,N10367);
not U3072 (N10550,N10354);
and U3073 (N10551,N10354,N3126);
nand U3074 (N10552,N7411,N10455);
and U3075 (N10553,N10375,N9539);
and U3076 (N10554,N10375,N9540);
and U3077 (N10555,N10375,N9541);
and U3078 (N10556,N10375,N6761);
not U3079 (N10557,N10406);
nand U3080 (N10558,N10406,N8243);
not U3081 (N10559,N10409);
nand U3082 (N10560,N10409,N8244);
not U3083 (N10561,N10412);
nand U3084 (N10562,N10412,N8245);
not U3085 (N10563,N10415);
nand U3086 (N10564,N10415,N8246);
nand U3087 (N10565,N7426,N10465);
not U3088 (N10566,N10419);
nand U3089 (N10567,N10419,N8248);
not U3090 (N10568,N10422);
nand U3091 (N10569,N10422,N8249);
not U3092 (N10570,N10425);
nand U3093 (N10571,N10425,N8250);
not U3094 (N10572,N10428);
nand U3095 (N10573,N10428,N8251);
not U3096 (N10574,N10399);
not U3097 (N10575,N10402);
not U3098 (N10576,N10388);
and U3099 (N10577,N10399,N10402,N10388);
and U3100 (N10581,N10360,N9543,N10273);
and U3101 (N10582,N10357,N9905,N10273);
not U3102 (N10583,N10367);
and U3103 (N10587,N10367,N5735);
and U3104 (N10588,N10367,N3135);
not U3105 (N10589,N10375);
and U3106 (N10594,N10381,N7180,N7159,N7170,N7149);
and U3107 (N10595,N10381,N7180,N7159,N7170);
and U3108 (N10596,N10381,N7180,N7170);
and U3109 (N10597,N10381,N7180);
and U3110 (N10598,N8444,N10381);
buff U3111 (N10602,N10381);
nand U3112 (N10609,N7479,N10515);
nand U3113 (N10610,N7491,N10517);
nand U3114 (N10621,N9149,N10534);
nand U3115 (N10626,N9206,N10542);
nand U3116 (N10627,N9223,N10544);
or U3117 (N10628,N10546,N10451);
and U3118 (N10629,N9733,N10547);
and U3119 (N10631,N5166,N10550);
nand U3120 (N10632,N10552,N10456);
nand U3121 (N10637,N7414,N10557);
nand U3122 (N10638,N7417,N10559);
nand U3123 (N10639,N7420,N10561);
nand U3124 (N10640,N7423,N10563);
nand U3125 (N10641,N10565,N10466);
nand U3126 (N10642,N7429,N10566);
nand U3127 (N10643,N7432,N10568);
nand U3128 (N10644,N7435,N10570);
nand U3129 (N10645,N7438,N10572);
and U3130 (N10647,N886,N887,N10577);
and U3131 (N10648,N10360,N8857,N10479);
and U3132 (N10649,N10357,N7609,N10479);
or U3133 (N10652,N8966,N10598);
or U3134 (N10659,N4675,N8451,N8452,N8453,N10594);
or U3135 (N10662,N4678,N8454,N8455,N10595);
or U3136 (N10665,N4682,N8456,N10596);
or U3137 (N10668,N4687,N10597);
not U3138 (N10671,N10509);
nand U3139 (N10672,N10509,N8615);
not U3140 (N10673,N10512);
nand U3141 (N10674,N10512,N8624);
nand U3142 (N10675,N10609,N10516);
nand U3143 (N10678,N10610,N10518);
not U3144 (N10681,N10519);
nand U3145 (N10682,N10519,N8644);
not U3146 (N10683,N10522);
nand U3147 (N10684,N10522,N8653);
not U3148 (N10685,N10525);
nand U3149 (N10686,N10525,N9454);
not U3150 (N10687,N10528);
nand U3151 (N10688,N10528,N9459);
not U3152 (N10689,N10531);
nand U3153 (N10690,N10531,N9978);
nand U3154 (N10691,N10621,N10535);
not U3155 (N10694,N10536);
nand U3156 (N10695,N10536,N9493);
not U3157 (N10696,N10539);
nand U3158 (N10697,N10539,N9498);
nand U3159 (N10698,N10626,N10543);
nand U3160 (N10701,N10627,N10545);
or U3161 (N10704,N10629,N10548);
and U3162 (N10705,N3159,N10583);
or U3163 (N10706,N10631,N10551);
and U3164 (N10707,N9737,N10589);
and U3165 (N10708,N9738,N10589);
and U3166 (N10709,N9243,N10589);
and U3167 (N10710,N5892,N10589);
nand U3168 (N10711,N10637,N10558);
nand U3169 (N10712,N10638,N10560);
nand U3170 (N10713,N10639,N10562);
nand U3171 (N10714,N10640,N10564);
nand U3172 (N10715,N10642,N10567);
nand U3173 (N10716,N10643,N10569);
nand U3174 (N10717,N10644,N10571);
nand U3175 (N10718,N10645,N10573);
not U3176 (N10719,N10602);
nand U3177 (N10720,N10602,N9244);
not U3178 (N10729,N10647);
and U3179 (N10730,N5178,N10583);
and U3180 (N10731,N2533,N10583);
nand U3181 (N10737,N7447,N10671);
nand U3182 (N10738,N7465,N10673);
or U3183 (N10739,N10648,N10649,N10581,N10582);
nand U3184 (N10746,N7503,N10681);
nand U3185 (N10747,N7521,N10683);
nand U3186 (N10748,N8678,N10685);
nand U3187 (N10749,N8690,N10687);
nand U3188 (N10750,N9685,N10689);
nand U3189 (N10753,N8757,N10694);
nand U3190 (N10754,N8769,N10696);
or U3191 (N10759,N10705,N10549);
or U3192 (N10760,N10707,N10553);
or U3193 (N10761,N10708,N10554);
or U3194 (N10762,N10709,N10555);
or U3195 (N10763,N10710,N10556);
nand U3196 (N10764,N8580,N10719);
and U3197 (N10765,N10652,N9890);
and U3198 (N10766,N10652,N9891);
and U3199 (N10767,N10652,N9892);
and U3200 (N10768,N10652,N8252);
not U3201 (N10769,N10659);
nand U3202 (N10770,N10659,N9245);
not U3203 (N10771,N10662);
nand U3204 (N10772,N10662,N9246);
not U3205 (N10773,N10665);
nand U3206 (N10774,N10665,N9247);
not U3207 (N10775,N10668);
nand U3208 (N10776,N10668,N9248);
or U3209 (N10778,N10730,N10587);
or U3210 (N10781,N10731,N10588);
not U3211 (N10784,N10652);
nand U3212 (N10789,N10737,N10672);
nand U3213 (N10792,N10738,N10674);
not U3214 (N10796,N10675);
nand U3215 (N10797,N10675,N8633);
not U3216 (N10798,N10678);
nand U3217 (N10799,N10678,N8638);
nand U3218 (N10800,N10746,N10682);
nand U3219 (N10803,N10747,N10684);
nand U3220 (N10806,N10748,N10686);
nand U3221 (N10809,N10749,N10688);
nand U3222 (N10812,N10750,N10690);
not U3223 (N10815,N10691);
nand U3224 (N10816,N10691,N9866);
nand U3225 (N10817,N10753,N10695);
nand U3226 (N10820,N10754,N10697);
not U3227 (N10823,N10698);
nand U3228 (N10824,N10698,N9505);
not U3229 (N10825,N10701);
nand U3230 (N10826,N10701,N9514);
nand U3231 (N10827,N10764,N10720);
nand U3232 (N10832,N8583,N10769);
nand U3233 (N10833,N8586,N10771);
nand U3234 (N10834,N8589,N10773);
nand U3235 (N10835,N8592,N10775);
not U3236 (N10836,N10739);
buff U3237 (N10837,N10778);
buff U3238 (N10838,N10778);
buff U3239 (N10839,N10781);
buff U3240 (N10840,N10781);
nand U3241 (N10845,N7482,N10796);
nand U3242 (N10846,N7494,N10798);
nand U3243 (N10857,N9473,N10815);
nand U3244 (N10862,N8781,N10823);
nand U3245 (N10863,N8799,N10825);
and U3246 (N10864,N10023,N10784);
and U3247 (N10865,N10024,N10784);
and U3248 (N10866,N9739,N10784);
and U3249 (N10867,N7136,N10784);
nand U3250 (N10868,N10832,N10770);
nand U3251 (N10869,N10833,N10772);
nand U3252 (N10870,N10834,N10774);
nand U3253 (N10871,N10835,N10776);
not U3254 (N10872,N10789);
nand U3255 (N10873,N10789,N8616);
not U3256 (N10874,N10792);
nand U3257 (N10875,N10792,N8625);
nand U3258 (N10876,N10845,N10797);
nand U3259 (N10879,N10846,N10799);
not U3260 (N10882,N10800);
nand U3261 (N10883,N10800,N8645);
not U3262 (N10884,N10803);
nand U3263 (N10885,N10803,N8654);
not U3264 (N10886,N10806);
nand U3265 (N10887,N10806,N9455);
not U3266 (N10888,N10809);
nand U3267 (N10889,N10809,N9460);
not U3268 (N10890,N10812);
nand U3269 (N10891,N10812,N9862);
nand U3270 (N10892,N10857,N10816);
not U3271 (N10895,N10817);
nand U3272 (N10896,N10817,N9494);
not U3273 (N10897,N10820);
nand U3274 (N10898,N10820,N9499);
nand U3275 (N10899,N10862,N10824);
nand U3276 (N10902,N10863,N10826);
or U3277 (N10905,N10864,N10765);
or U3278 (N10906,N10865,N10766);
or U3279 (N10907,N10866,N10767);
or U3280 (N10908,N10867,N10768);
nand U3281 (N10909,N7450,N10872);
nand U3282 (N10910,N7468,N10874);
nand U3283 (N10915,N7506,N10882);
nand U3284 (N10916,N7524,N10884);
nand U3285 (N10917,N8681,N10886);
nand U3286 (N10918,N8693,N10888);
nand U3287 (N10919,N9462,N10890);
nand U3288 (N10922,N8760,N10895);
nand U3289 (N10923,N8772,N10897);
nand U3290 (N10928,N10909,N10873);
nand U3291 (N10931,N10910,N10875);
not U3292 (N10934,N10876);
nand U3293 (N10935,N10876,N8634);
not U3294 (N10936,N10879);
nand U3295 (N10937,N10879,N8639);
nand U3296 (N10938,N10915,N10883);
nand U3297 (N10941,N10916,N10885);
nand U3298 (N10944,N10917,N10887);
nand U3299 (N10947,N10918,N10889);
nand U3300 (N10950,N10919,N10891);
not U3301 (N10953,N10892);
nand U3302 (N10954,N10892,N9476);
nand U3303 (N10955,N10922,N10896);
nand U3304 (N10958,N10923,N10898);
not U3305 (N10961,N10899);
nand U3306 (N10962,N10899,N9506);
not U3307 (N10963,N10902);
nand U3308 (N10964,N10902,N9515);
nand U3309 (N10969,N7485,N10934);
nand U3310 (N10970,N7497,N10936);
nand U3311 (N10981,N8718,N10953);
nand U3312 (N10986,N8784,N10961);
nand U3313 (N10987,N8802,N10963);
not U3314 (N10988,N10928);
nand U3315 (N10989,N10928,N8617);
not U3316 (N10990,N10931);
nand U3317 (N10991,N10931,N8626);
nand U3318 (N10992,N10969,N10935);
nand U3319 (N10995,N10970,N10937);
not U3320 (N10998,N10938);
nand U3321 (N10999,N10938,N8646);
not U3322 (N11000,N10941);
nand U3323 (N11001,N10941,N8655);
not U3324 (N11002,N10944);
nand U3325 (N11003,N10944,N9456);
not U3326 (N11004,N10947);
nand U3327 (N11005,N10947,N9461);
not U3328 (N11006,N10950);
nand U3329 (N11007,N10950,N9465);
nand U3330 (N11008,N10981,N10954);
not U3331 (N11011,N10955);
nand U3332 (N11012,N10955,N9495);
not U3333 (N11013,N10958);
nand U3334 (N11014,N10958,N9500);
nand U3335 (N11015,N10986,N10962);
nand U3336 (N11018,N10987,N10964);
nand U3337 (N11023,N7453,N10988);
nand U3338 (N11024,N7471,N10990);
nand U3339 (N11027,N7509,N10998);
nand U3340 (N11028,N7527,N11000);
nand U3341 (N11029,N8684,N11002);
nand U3342 (N11030,N8696,N11004);
nand U3343 (N11031,N8702,N11006);
nand U3344 (N11034,N8763,N11011);
nand U3345 (N11035,N8775,N11013);
not U3346 (N11040,N10992);
nand U3347 (N11041,N10992,N8294);
not U3348 (N11042,N10995);
nand U3349 (N11043,N10995,N8295);
nand U3350 (N11044,N11023,N10989);
nand U3351 (N11047,N11024,N10991);
nand U3352 (N11050,N11027,N10999);
nand U3353 (N11053,N11028,N11001);
nand U3354 (N11056,N11029,N11003);
nand U3355 (N11059,N11030,N11005);
nand U3356 (N11062,N11031,N11007);
not U3357 (N11065,N11008);
nand U3358 (N11066,N11008,N9477);
nand U3359 (N11067,N11034,N11012);
nand U3360 (N11070,N11035,N11014);
not U3361 (N11073,N11015);
nand U3362 (N11074,N11015,N9507);
not U3363 (N11075,N11018);
nand U3364 (N11076,N11018,N9516);
nand U3365 (N11077,N7488,N11040);
nand U3366 (N11078,N7500,N11042);
nand U3367 (N11095,N8721,N11065);
nand U3368 (N11098,N8787,N11073);
nand U3369 (N11099,N8805,N11075);
nand U3370 (N11100,N11077,N11041);
nand U3371 (N11103,N11078,N11043);
not U3372 (N11106,N11056);
nand U3373 (N11107,N11056,N9319);
not U3374 (N11108,N11059);
nand U3375 (N11109,N11059,N9320);
not U3376 (N11110,N11067);
nand U3377 (N11111,N11067,N9381);
not U3378 (N11112,N11070);
nand U3379 (N11113,N11070,N9382);
not U3380 (N11114,N11044);
nand U3381 (N11115,N11044,N8618);
not U3382 (N11116,N11047);
nand U3383 (N11117,N11047,N8619);
not U3384 (N11118,N11050);
nand U3385 (N11119,N11050,N8647);
not U3386 (N11120,N11053);
nand U3387 (N11121,N11053,N8648);
not U3388 (N11122,N11062);
nand U3389 (N11123,N11062,N9466);
nand U3390 (N11124,N11095,N11066);
nand U3391 (N11127,N11098,N11074);
nand U3392 (N11130,N11099,N11076);
nand U3393 (N11137,N8687,N11106);
nand U3394 (N11138,N8699,N11108);
nand U3395 (N11139,N8766,N11110);
nand U3396 (N11140,N8778,N11112);
nand U3397 (N11141,N7456,N11114);
nand U3398 (N11142,N7474,N11116);
nand U3399 (N11143,N7512,N11118);
nand U3400 (N11144,N7530,N11120);
nand U3401 (N11145,N8705,N11122);
and U3402 (N11152,N11103,N8871,N10283);
and U3403 (N11153,N11100,N7655,N10283);
and U3404 (N11154,N11103,N9551,N10119);
and U3405 (N11155,N11100,N9917,N10119);
nand U3406 (N11156,N11137,N11107);
nand U3407 (N11159,N11138,N11109);
nand U3408 (N11162,N11139,N11111);
nand U3409 (N11165,N11140,N11113);
nand U3410 (N11168,N11141,N11115);
nand U3411 (N11171,N11142,N11117);
nand U3412 (N11174,N11143,N11119);
nand U3413 (N11177,N11144,N11121);
nand U3414 (N11180,N11145,N11123);
not U3415 (N11183,N11124);
nand U3416 (N11184,N11124,N9468);
not U3417 (N11185,N11127);
nand U3418 (N11186,N11127,N9508);
not U3419 (N11187,N11130);
nand U3420 (N11188,N11130,N9509);
or U3421 (N11205,N11152,N11153,N11154,N11155);
nand U3422 (N11210,N8724,N11183);
nand U3423 (N11211,N8790,N11185);
nand U3424 (N11212,N8808,N11187);
not U3425 (N11213,N11168);
nand U3426 (N11214,N11168,N8260);
not U3427 (N11215,N11171);
nand U3428 (N11216,N11171,N8261);
not U3429 (N11217,N11174);
nand U3430 (N11218,N11174,N8296);
not U3431 (N11219,N11177);
nand U3432 (N11220,N11177,N8297);
and U3433 (N11222,N11159,N9575,N1218);
and U3434 (N11223,N11156,N8927,N1218);
and U3435 (N11224,N11159,N9935,N750);
and U3436 (N11225,N11156,N10132,N750);
and U3437 (N11226,N11165,N9608,N10497);
and U3438 (N11227,N11162,N9001,N10497);
and U3439 (N11228,N11165,N9949,N10301);
and U3440 (N11229,N11162,N10160,N10301);
not U3441 (N11231,N11180);
nand U3442 (N11232,N11180,N9467);
nand U3443 (N11233,N11210,N11184);
nand U3444 (N11236,N11211,N11186);
nand U3445 (N11239,N11212,N11188);
nand U3446 (N11242,N7459,N11213);
nand U3447 (N11243,N7462,N11215);
nand U3448 (N11244,N7515,N11217);
nand U3449 (N11245,N7518,N11219);
not U3450 (N11246,N11205);
nand U3451 (N11250,N8708,N11231);
or U3452 (N11252,N11222,N11223,N11224,N11225);
or U3453 (N11257,N11226,N11227,N11228,N11229);
nand U3454 (N11260,N11242,N11214);
nand U3455 (N11261,N11243,N11216);
nand U3456 (N11262,N11244,N11218);
nand U3457 (N11263,N11245,N11220);
not U3458 (N11264,N11233);
nand U3459 (N11265,N11233,N9322);
not U3460 (N11267,N11236);
nand U3461 (N11268,N11236,N9383);
not U3462 (N11269,N11239);
nand U3463 (N11270,N11239,N9384);
nand U3464 (N11272,N11250,N11232);
not U3465 (N11277,N11261);
and U3466 (N11278,N10273,N11260);
not U3467 (N11279,N11263);
and U3468 (N11280,N10119,N11262);
nand U3469 (N11282,N8714,N11264);
not U3470 (N11283,N11252);
nand U3471 (N11284,N8793,N11267);
nand U3472 (N11285,N8796,N11269);
not U3473 (N11286,N11257);
and U3474 (N11288,N11277,N10479);
and U3475 (N11289,N11279,N10283);
not U3476 (N11290,N11272);
nand U3477 (N11291,N11272,N9321);
nand U3478 (N11292,N11282,N11265);
nand U3479 (N11293,N11284,N11268);
nand U3480 (N11294,N11285,N11270);
nand U3481 (N11295,N8711,N11290);
not U3482 (N11296,N11292);
not U3483 (N11297,N11294);
and U3484 (N11298,N10301,N11293);
or U3485 (N11299,N11288,N11278);
or U3486 (N11302,N11289,N11280);
nand U3487 (N11307,N11295,N11291);
and U3488 (N11308,N11296,N1218);
and U3489 (N11309,N11297,N10497);
nand U3490 (N11312,N11302,N11246);
nand U3491 (N11313,N11299,N10836);
not U3492 (N11314,N11299);
not U3493 (N11315,N11302);
and U3494 (N11316,N750,N11307);
or U3495 (N11317,N11309,N11298);
nand U3496 (N11320,N11205,N11315);
nand U3497 (N11321,N10739,N11314);
or U3498 (N11323,N11308,N11316);
nand U3499 (N11327,N11312,N11320);
nand U3500 (N11328,N11313,N11321);
nand U3501 (N11329,N11317,N11286);
not U3502 (N11331,N11317);
not U3503 (N11333,N11327);
not U3504 (N11334,N11328);
nand U3505 (N11335,N11257,N11331);
nand U3506 (N11336,N11323,N11283);
not U3507 (N11337,N11323);
nand U3508 (N11338,N11329,N11335);
nand U3509 (N11339,N11252,N11337);
not U3510 (N11340,N11338);
nand U3511 (N11341,N11336,N11339);
not U3512 (N11342,N11341);
buff U3513 (B241,N241);
endmodule
