module c2670 ( N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N138, N139, N140, N141, N142, N219, N224, N227, N230, N231, N234, N237, N241, N246, N253, N256, N259, N262, N263, N266, N269, N272, N275, N278, N281, N284, N287, N290, N294, N297, N301, N305, N309, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N143_I, N144_I, N145_I, N146_I, N147_I, N148_I, N149_I, N150_I, N151_I, N152_I, N153_I, N154_I, N155_I, N156_I, N157_I, N158_I, N159_I, N160_I, N161_I, N162_I, N163_I, N164_I, N165_I, N166_I, N167_I, N168_I, N169_I, N170_I, N171_I, N172_I, N173_I, N174_I, N175_I, N176_I, N177_I, N178_I, N179_I, N180_I, N181_I, N182_I, N183_I, N184_I, N185_I, N186_I, N187_I, N188_I, N189_I, N190_I, N191_I, N192_I, N193_I, N194_I, N195_I, N196_I, N197_I, N198_I, N199_I, N200_I, N201_I, N202_I, N203_I, N204_I, N205_I, N206_I, N207_I, N208_I, N209_I, N210_I, N211_I, N212_I, N213_I, N214_I, N215_I, N216_I, N217_I, N218_I, N398, N400, N401, N419, N420, N456, N457, N458, N487, N488, N489, N490, N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029, N1269, N1277, N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821, N1969, N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022, N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, N2970, N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3881, N3882, N143_O, N144_O, N145_O, N146_O, N147_O, N148_O, N149_O, N150_O, N151_O, N152_O, N153_O, N154_O, N155_O, N156_O, N157_O, N158_O, N159_O, N160_O, N161_O, N162_O, N163_O, N164_O, N165_O, N166_O, N167_O, N168_O, N169_O, N170_O, N171_O, N172_O, N173_O, N174_O, N175_O, N176_O, N177_O, N178_O, N179_O, N180_O, N181_O, N182_O, N183_O, N184_O, N185_O, N186_O, N187_O, N188_O, N189_O, N190_O, N191_O, N192_O, N193_O, N194_O, N195_O, N196_O, N197_O, N198_O, N199_O, N200_O, N201_O, N202_O, N203_O, N204_O, N205_O, N206_O, N207_O, N208_O, N209_O, N210_O, N211_O, N212_O, N213_O, N214_O, N215_O, N216_O, N217_O, N218_O);
input N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,N216_I,N217_I,N218_I;
output N398,N400,N401,N419,N420,N456,N457,N458,N487,N488,N489,N490,N491,N492,N493,N494,N792,N799,N805,N1026,N1028,N1029,N1269,N1277,N1448,N1726,N1816,N1817,N1818,N1819,N1820,N1821,N1969,N1970,N1971,N2010,N2012,N2014,N2016,N2018,N2020,N2022,N2387,N2388,N2389,N2390,N2496,N2643,N2644,N2891,N2925,N2970,N2971,N3038,N3079,N3546,N3671,N3803,N3804,N3809,N3851,N3881,N3882,N143_O,N144_O,N145_O,N146_O,N147_O,N148_O,N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,N156_O,N157_O,N158_O,N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,N166_O,N167_O,N168_O,N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,N176_O,N177_O,N178_O,N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,N186_O,N187_O,N188_O,N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,N196_O,N197_O,N198_O,N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,N206_O,N207_O,N208_O,N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,N216_O,N217_O,N218_O;
wire n279,n280,n281,n282,n283,n284,n285,n286,n288,n289,n290,n291,n292,n293,n294,n295,n296,n297,n298,n299,n300,n301,n302,n303,n304,n305,n306,n307,n308,n309,n310,n311,n312,n313,n314,n315,n316,n317,n318,n319,n320,n321,n322,n323,n324,n325,n326,n327,n328,n329,n330,n331,n332,n333,n334,n335,n336,n337,n338,n339,n340,n341,n342,n343,n344,n345,n346,n347,n348,n349,n350,n351,n352,n353,n354,n355,n356,n357,n358,n359,n360,n361,n362,n363,n364,n365,n366,n367,n368,n369,n370,n371,n372,n373,n374,n375,n376,n377,n378,n379,n380,n381,n382,n383,n384,n385,n386,n387,n388,n389,n390,n391,n392,n393,n394,n395,n396,n397,n398,n399,n400,n401,n402,n403,n404,n405,n406,n407,n408,n409,n410,n411,n412,n413,n414,n415,n416,n417,n418,n419,n420,n421,n422,n423,n424,n425,n426,n427,n428,n429,n430,n431,n432,n433,n434,n435,n436,n437,n438,n439,n440,n441,n442,n443,n444,n445,n446,n447,n448,n449,n450,n451,n452,n453,n454,n455,n456,n457,n458,n459,n460,n461,n462,n463,n464,n465,n466,n467,n468,n469,n470,n471,n472,n473,n474,n475,n476,n477,n478,n479,n480,n481,n482,n483,n484,n485,n486,n487,n488,n489,n490,n491,n492,n493,n494,n495,n496,n497,n498,n499,n500,n501,n502,n503,n504,n505,n506,n507,n508,n509,n510,n511,n512,n513,n514,n515,n516,n517,n518,n519,n520,n521,n522,n523,n524,n525,n526,n527,n528,n529,n530,n531,n532,n533,n534,n535,n536,n537,n538,n539,n540,n541,n542,n543,n544,n545,n546,n547,n548,n549,n550,n551,n552,n553,n554,n555,n556,n557,n558,n559,n560,n561,n562,n563,n564,n565,n566,n567,n568,n569,n570,n571,n572,n573,n574,n575,n576,n577,n578,n579,n580,n581,n582,n583,n584,n585,n586,n587,n588,n589,n590,n591,n592,n593,n594,n595,n596,n597,n598,n599,n600,n601,n602,n603,n604,n605,n606,n607,n608,n609,n610,n611,n612,n613,n614,n615,n616,n617,n618,n619,n620,n621,n622,n623,n624,n625,n626,n627,n628,n629,n630,n631,n632,n633,n634,n635,n636,n637,n638,n639,n640,n641,n642,n643,n644,n645,n646,n647,n648,n649,n650,n651,n652,n653,n654,n655,n656,n657,n658,n659,n660,n661,n662,n663,n664,n665,n666,n667,n668,n669,n670,n671,n672,n673,n674,n675,n676,n677,n678,n679,n680,n681,n682,n683,n684,n685,n686,n687,n688,n689,n690,n691,n692,n693,n694,n695,n696,n697,n698,n699,n700,n701,n702,n703,n704,n705,n706,n707,n708,n709,n710,n711,n712,n713,n714,n715,n716,n717,n718,n719,n720,n721,n722,n723,n724,n725,n726,n727,n728,n729,n730,n731,n732,n733,n734,n735,n736,n737,n738,n739,n740,n741,n742,n743,n744,n745,n746,n747,n748,n749,n750,n751,n752,n753,n754,n755,n756,n757,n758,n759,n760,n761,n762,n763,n764,n765,n766,n767,n768,n769,n770,n771,n772,n773,n774,n775,n776,n777,n778,n779,n780,n781,n782,n783,n784,n785,n786,n787,n788,n789,n790,n791,n792,n793,n794,n795,n796,n797,n798,n799,n800,n801,n802,n803,n804,n805,n806,n807,n808,n809,n810,n811,n812,n813,n814,n815,n816,n817,n818,n819,n820,n821,n822,n823,n824,n825,n826,n827,n828,n829,n830,n831,n832,n833,n834,n835,n836,n837,n838,n839,n840,n841,n842,n843,n844,n845,n846,n847,n848,n849,n850,n851,n852,n853,n854,n855,n856,n857,n858,n859,n860,n861,n862,n863,n864,n865,n866,n867,n868,n869,n870,n871,n872,n873,n874,n875,n876,n877,n878,n879,n880,n881,n882,n883,n884,n885,n886,n887,n888,n889,n890,n891,n892,n893,n894,n895,n896,n897,n898,n899,n900,n901,n902,n903,n904,n905,n906,n907,n908,n909,n910,n911,n912,n913,n914,n915;
  
buff U688 (N398, N219);
buff U689 (N400, N219);
buff U690 (N401, N219);
buff U691 (N419, N253);
buff U692 (N420, N253);
buff U693 (N456, N290);
buff U694 (N457, N290);
buff U695 (N458, N290);
buff U696 (N805, N219);
buff U697 (N2388, N2387);
buff U698 (N2390, N2389);
buff U699 (N2644, N2643);
buff U700 (N3804, N3803);
buff U701 (N143_O, N143_I);
buff U702 (N144_O, N144_I);
buff U703 (N145_O, N145_I);
buff U704 (N146_O, N146_I);
buff U705 (N147_O, N147_I);
buff U706 (N148_O, N148_I);
buff U707 (N149_O, N149_I);
buff U708 (N150_O, N150_I);
buff U709 (N151_O, N151_I);
buff U710 (N152_O, N152_I);
buff U711 (N153_O, N153_I);
buff U712 (N154_O, N154_I);
buff U713 (N155_O, N155_I);
buff U714 (N156_O, N156_I);
buff U715 (N157_O, N157_I);
buff U716 (N158_O, N158_I);
buff U717 (N159_O, N159_I);
buff U718 (N160_O, N160_I);
buff U719 (N161_O, N161_I);
buff U720 (N162_O, N162_I);
buff U721 (N163_O, N163_I);
buff U722 (N164_O, N164_I);
buff U723 (N165_O, N165_I);
buff U724 (N166_O, N166_I);
buff U725 (N167_O, N167_I);
buff U726 (N168_O, N168_I);
buff U727 (N169_O, N169_I);
buff U728 (N170_O, N170_I);
buff U729 (N171_O, N171_I);
buff U730 (N172_O, N172_I);
buff U731 (N173_O, N173_I);
buff U732 (N174_O, N174_I);
buff U733 (N175_O, N175_I);
buff U734 (N176_O, N176_I);
buff U735 (N177_O, N177_I);
buff U736 (N178_O, N178_I);
buff U737 (N179_O, N179_I);
buff U738 (N180_O, N180_I);
buff U739 (N181_O, N181_I);
buff U740 (N182_O, N182_I);
buff U741 (N183_O, N183_I);
buff U742 (N184_O, N184_I);
buff U743 (N185_O, N185_I);
buff U744 (N186_O, N186_I);
buff U745 (N187_O, N187_I);
buff U746 (N188_O, N188_I);
buff U747 (N189_O, N189_I);
buff U748 (N190_O, N190_I);
buff U749 (N191_O, N191_I);
buff U750 (N192_O, N192_I);
buff U751 (N193_O, N193_I);
buff U752 (N194_O, N194_I);
buff U753 (N195_O, N195_I);
buff U754 (N196_O, N196_I);
buff U755 (N197_O, N197_I);
buff U756 (N198_O, N198_I);
buff U757 (N199_O, N199_I);
buff U758 (N200_O, N200_I);
buff U759 (N201_O, N201_I);
buff U760 (N202_O, N202_I);
buff U761 (N203_O, N203_I);
buff U762 (N204_O, N204_I);
buff U763 (N205_O, N205_I);
buff U764 (N206_O, N206_I);
buff U765 (N207_O, N207_I);
buff U766 (N208_O, N208_I);
buff U767 (N209_O, N209_I);
buff U768 (N210_O, N210_I);
buff U769 (N211_O, N211_I);
buff U770 (N212_O, N212_I);
buff U771 (N213_O, N213_I);
buff U772 (N214_O, N214_I);
buff U773 (N215_O, N215_I);
buff U774 (N216_O, N216_I);
buff U775 (N217_O, N217_I);
buff U776 (N218_O, N218_I);
nor U1 (N3038, n279, n280);
not U2 (N2022, n281);
not U3 (N2020, n282);
not U4 (N2018, n283);
not U5 (N2016, N1819);
not U6 (N2014, N1820);
not U7 (N2012, N1821);
not U8 (N2010, n284);
nor U9 (N3881, n285, n286);
nand U11 (N3851, n288, n289);
not U12 (N3079, N3038);
nand U13 (N2891, n290, n291);
nand U14 (N1971, n292, n293);
nand U15 (N1970, N36, n292);
nand U16 (N1969, N241, n294);
nor U17 (N1277, n295, n296);
nand U18 (N1029, N231, n297);
nand U19 (N1269, N325, n297);
nand U20 (N792, n298, n299);
nand U21 (N1028, N7, N237);
not U22 (N494, N108);
not U23 (N493, N57);
not U24 (N492, N120);
not U25 (N491, N69);
not U26 (N490, N96);
not U27 (N489, N82);
not U28 (N488, N132);
not U29 (N487, N44);
nand U30 (N799, N237, n300);
nor U31 (n301, n302, n303);
nor U32 (N1816, n304, n305);
nor U33 (N1817, n306, n307);
nor U34 (n308, n309, n310);
nor U35 (n311, n312, n313);
nor U36 (n314, n315, n316);
nor U37 (n317, n318, n319);
nor U38 (n320, n321, n322);
nor U39 (N1818, n323, n324);
nor U40 (N1820, n325, n326);
nor U41 (N1821, n327, n328);
nor U42 (n329, n330, n331);
nor U43 (n294, n332, n333);
nor U44 (n284, n334, n335);
nor U45 (n336, n337, n338);
nor U46 (n281, n339, n340);
nor U47 (n282, n341, n342);
nor U48 (n283, n343, n344);
nor U49 (N1819, n345, n346);
nor U50 (n347, N262, N1818);
nor U51 (n348, n349, n350);
nor U52 (n351, n352, n353);
nor U53 (n354, n352, n355);
nor U54 (n356, n357, n358);
nand U55 (n359, n360, n361);
nor U56 (n362, N1821, n363);
nand U57 (n364, n365, n366);
nor U58 (n367, n368, n369);
nor U59 (n370, n371, n372);
nor U60 (n373, n367, n370);
nor U61 (n374, n352, n375);
nor U62 (n376, n354, n373);
nor U63 (n377, n374, n376);
nor U64 (n378, n352, n379);
nor U65 (n380, n351, n377);
nor U66 (n381, n378, n380);
nor U67 (n382, n383, n384);
nor U68 (n385, n386, n387);
nor U69 (n388, n389, n390);
nor U70 (n391, n392, n393);
nor U71 (n394, n395, n396);
nand U72 (N2496, n336, n397);
nor U73 (n398, n284, n359);
nor U74 (n371, n356, n394);
not U75 (n399, n336);
not U76 (n400, N301);
not U77 (n401, N297);
not U78 (n402, N309);
not U79 (n403, N305);
nor U80 (n404, N319, N322);
not U81 (n405, N319);
nor U82 (n406, n405, N322);
nor U83 (n407, n408, N319);
nor U84 (n409, n408, n405);
not U85 (n410, n314);
not U86 (n411, n317);
not U87 (n412, N1816);
not U88 (n413, n308);
nor U89 (n414, N227, N234);
not U90 (n415, N227);
nor U91 (n416, n417, n415);
nor U92 (n418, n415, N234);
nor U93 (n419, n417, N227);
not U94 (n420, n329);
not U95 (n421, n294);
not U96 (n422, N294);
not U97 (n423, N275);
not U98 (n424, N266);
not U99 (n425, N284);
not U100 (n426, N287);
not U101 (n427, N278);
not U102 (n428, N281);
not U103 (n429, N263);
nand U104 (n430, n431, n432);
nand U105 (n349, n433, N40);
not U106 (n357, N8);
nand U107 (n352, N8, n434);
nand U108 (n369, n435, N8);
nor U109 (n368, n357, N1819);
nand U110 (n436, n437, n294);
nor U111 (n395, n357, N1820);
nor U112 (n438, n399, N230);
nor U113 (n292, n439, n440);
not U114 (n441, N241);
nand U115 (n296, n442, n443);
nand U116 (n295, n444, n445);
nor U117 (n446, n447, n448);
nor U118 (n449, n450, n451);
nand U119 (N2971, n452, n453);
nand U120 (n454, n455, n456);
nand U121 (n457, n458, n459);
nand U122 (n460, n461, n462);
nand U123 (n463, n464, n465);
nand U124 (n466, n467, n468);
nand U125 (n469, n470, n471);
nand U126 (n472, n473, n474);
nand U127 (n475, n476, n477);
nand U128 (n478, n375, n355);
nand U129 (n479, n480, n481);
nand U130 (n482, n483, n350);
nand U131 (n484, n379, n353);
nand U132 (n363, n485, n486);
nand U133 (n358, n487, n488);
nand U134 (N3803, n489, n490);
nand U135 (n491, n492, n493);
nand U136 (N2643, n494, n495);
nand U137 (N2389, n496, n497);
nand U138 (N2387, n498, n499);
nand U139 (n500, N2, N15);
nor U140 (n299, n400, n401);
nor U141 (n298, n402, n403);
nand U142 (n312, n501, n502);
nand U143 (n313, n503, n504);
nand U144 (n315, n505, n506);
nand U145 (n316, n507, n508);
nand U146 (n318, n509, n510);
nand U147 (n319, n511, n512);
nand U148 (n302, n513, n514);
nand U149 (n303, n515, n516);
nand U150 (n304, n517, n518);
nand U151 (n305, n519, n520);
nand U152 (n306, n521, n522);
nand U153 (n307, n523, n524);
nand U154 (n309, n525, n526);
nand U155 (n310, n527, n528);
nand U156 (n321, n529, n530);
nand U157 (n322, n531, n532);
nand U158 (n323, n533, n534);
nand U159 (n324, n535, n536);
nand U160 (n537, n538, n539);
nor U161 (n540, n541, n542);
nand U162 (n543, n544, n545);
nor U163 (n546, n547, n548);
nor U164 (n549, n550, n551);
nand U165 (n552, n553, n554);
nand U166 (n325, n555, n556);
nand U167 (n326, n557, n558);
nand U168 (n327, n559, n560);
nand U169 (n328, n561, n562);
nand U170 (n339, n563, n564);
nand U171 (n340, n565, n566);
nand U172 (n341, n567, n568);
nand U173 (n342, n569, n570);
nand U174 (n343, n571, n572);
nand U175 (n344, n573, n574);
nand U176 (n345, n575, n576);
nand U177 (n346, n577, n578);
nand U178 (n330, n579, n580);
nand U179 (n331, n581, n582);
nand U180 (n332, n583, n584);
nand U181 (n333, n585, n586);
nand U182 (n334, n587, n588);
nand U183 (n335, n589, n590);
nand U184 (n337, n591, n592);
nand U185 (n338, n593, n594);
nand U186 (n595, n596, n597);
nand U187 (n598, n599, n600);
nand U188 (n601, n602, n603);
nor U189 (n604, n605, n606);
nand U190 (n607, n608, n609);
nor U191 (n610, n611, n612);
nor U192 (n613, n614, n615);
nand U193 (n616, n617, n618);
nand U194 (n619, n620, n621);
nand U195 (n622, n623, n624);
nand U196 (n625, n626, n627);
nor U197 (n628, n629, n630);
nand U198 (n631, n632, n633);
nand U199 (n634, n635, n636);
nand U200 (n637, n638, n639);
nand U201 (n640, n641, n642);
nand U202 (n643, n644, n645);
nand U203 (n646, n647, n648);
nor U204 (n649, n650, n651);
nor U205 (n652, n653, n654);
nor U206 (n443, N490, N489);
nor U207 (n442, N488, N487);
nor U208 (n445, N494, N493);
nor U209 (n444, N492, N491);
nor U210 (n655, N3809, N3671);
nand U211 (n286, n656, n655);
nor U212 (n657, N2971, N2970);
nand U213 (n285, N1726, n657);
nor U214 (n433, n347, n412);
nor U215 (n658, N294, n411);
nor U216 (n659, n317, n422);
nor U217 (n660, n314, n426);
nor U218 (n661, n308, n425);
nand U219 (n662, N1816, N40);
nor U220 (n663, n362, n398);
nand U221 (n372, n664, n665);
nand U222 (n666, n667, n668);
nor U223 (n669, n348, n381);
nor U224 (n670, N2022, N281);
nand U225 (n671, n672, n673);
nand U226 (n674, n675, n676);
nor U227 (n677, n678, n679);
nor U228 (n680, n681, n682);
nand U229 (n386, n680, n677);
nor U230 (n683, n684, n685);
nand U231 (n387, n683, N28);
nor U232 (n686, n301, n454);
nor U233 (n687, n457, n460);
nand U234 (n383, n687, n686);
nor U235 (n688, n463, n466);
nand U236 (n384, n688, n689);
nand U237 (n690, n691, n692);
nor U238 (n693, n694, n690);
nor U239 (n695, n696, n697);
nand U240 (n392, n695, n693);
nor U241 (n698, n699, n700);
nor U242 (n701, n702, n703);
nand U243 (n393, n701, n698);
nand U244 (n704, n705, n706);
nor U245 (n707, n469, n704);
nor U246 (n708, n472, n475);
nand U247 (n389, n708, n707);
nor U248 (n709, n478, n479);
nor U249 (n710, n482, n484);
nand U250 (n390, n710, n709);
nand U251 (n279, n711, N11);
nand U252 (n280, n712, n713);
nand U253 (n439, N237, N1726);
not U254 (n714, N256);
not U255 (n715, N259);
not U256 (n716, N346);
not U257 (n717, N349);
nor U258 (n718, N349, n716);
nor U259 (n719, N346, n717);
nor U260 (n720, n718, n719);
nor U261 (n721, N259, n714);
nor U262 (n722, N256, n715);
nor U263 (n723, n721, n722);
nand U264 (n724, n725, n726);
not U265 (n727, n301);
not U266 (n728, N1817);
not U267 (n729, n320);
not U268 (n730, N1818);
nor U269 (n731, n552, n549);
nand U270 (n732, n549, n552);
nand U271 (n733, n734, n732);
nor U272 (n735, N2018, N1819);
nor U273 (n736, N2016, n283);
nor U274 (n737, n735, n736);
nor U275 (n738, N2022, n282);
nor U276 (n739, N2020, n281);
nor U277 (n740, n738, n739);
nand U278 (n741, n742, n743);
not U279 (n744, N313);
not U280 (n291, N316);
not U281 (n745, N272);
not U282 (n746, N269);
nor U283 (n747, N281, n427);
nor U284 (n748, N278, n428);
nor U285 (n749, n747, n748);
nor U286 (n750, N287, n425);
nor U287 (n751, N284, n426);
nor U288 (n752, n750, n751);
nand U289 (n753, n754, n755);
nor U290 (n756, n662, n757);
nor U291 (n758, n756, n745);
nor U292 (n759, n402, n434);
nor U293 (n435, n758, n759);
nor U294 (n760, n756, n714);
nor U295 (n761, n426, n434);
nor U296 (n437, n760, n761);
nor U297 (n762, n756, n715);
nor U298 (n763, n422, n434);
nor U299 (n764, n762, n763);
nor U300 (n765, N297, n434);
nor U301 (n766, n756, N263);
nor U302 (n767, n765, n766);
not U303 (n768, N246);
nand U304 (n769, n770, n441);
nor U305 (n771, n772, n420);
nor U306 (n773, n329, n769);
nor U307 (N3546, n771, n773);
not U308 (n774, N29);
nor U309 (n775, N32, n426);
nor U310 (n776, N287, n777);
nor U311 (n678, n775, n776);
nor U312 (n778, N26, n422);
nor U313 (n779, N294, n780);
nor U314 (n679, n778, n779);
nor U315 (n781, N33, n401);
nor U316 (n782, N297, n783);
nor U317 (n681, n781, n782);
nor U318 (n784, N35, n402);
nor U319 (n785, N309, n786);
nor U320 (n682, n784, n785);
nor U321 (n787, N27, n400);
nor U322 (n788, N301, n789);
nor U323 (n684, n787, n788);
nor U324 (n790, N34, n403);
nor U325 (n791, N305, n792);
nor U326 (n685, n790, n791);
nor U327 (n793, N1817, n402);
nor U328 (n794, N309, n728);
nor U329 (n689, n793, n794);
nor U330 (n795, n382, n774);
nor U331 (n796, N29, n385);
nor U332 (n713, n795, n796);
nor U333 (n797, N4, n715);
nor U334 (n798, N259, n799);
nor U335 (n694, n797, n798);
nor U336 (n800, N5, n424);
nor U337 (n801, N266, n802);
nor U338 (n696, n800, n801);
nor U339 (n803, N21, n746);
nor U340 (n804, N269, n805);
nor U341 (n697, n803, n804);
nor U342 (n806, N22, n745);
nor U343 (n807, N272, n808);
nor U344 (n699, n806, n807);
nor U345 (n809, N23, n423);
nor U346 (n810, N275, n811);
nor U347 (n700, n809, n810);
nor U348 (n812, N6, n427);
nor U349 (n813, N278, n814);
nor U350 (n702, n812, n813);
nor U351 (n815, N24, n428);
nor U352 (n816, N281, n817);
nor U353 (n703, n815, n816);
nor U354 (n818, n284, n429);
nor U355 (n819, N2010, N263);
nor U356 (n706, n818, n819);
nor U357 (n820, n336, n715);
nor U358 (n821, N259, n399);
nor U359 (n705, n820, n821);
not U360 (n822, N16);
nor U361 (n823, n388, n822);
nor U362 (n824, N16, n391);
nor U363 (n712, n823, n824);
nor U364 (n825, n301, n744);
nor U365 (n826, N313, n727);
nor U366 (n290, n825, n826);
not U367 (N3882, N3881);
not U368 (n434, n756);
nand U369 (n827, N219, N94);
not U370 (N1026, n827);
not U371 (n572, n419);
nand U372 (n514, N135, n404);
nand U373 (n513, N99, n406);
nand U374 (n516, N123, n407);
nand U375 (n515, N111, n409);
nand U376 (n518, N137, n404);
nand U377 (n517, N101, n406);
nand U378 (n520, N125, n407);
nand U379 (n519, N113, n409);
nand U380 (n522, N136, n404);
nand U381 (n521, N100, n406);
nand U382 (n524, N124, n407);
nand U383 (n523, N112, n409);
nand U384 (n526, N131, n404);
nand U385 (n525, N95, n406);
nand U386 (n528, N119, n407);
nand U387 (n527, N107, n409);
nand U388 (n502, N142, n404);
nand U389 (n501, N106, n406);
nand U390 (n504, N130, n407);
nand U391 (n503, N118, n409);
nand U392 (n506, N141, n404);
nand U393 (n505, N105, n406);
nand U394 (n508, N129, n407);
nand U395 (n507, N117, n409);
nand U396 (n510, N140, n404);
nand U397 (n509, N104, n406);
nand U398 (n512, N128, n407);
nand U399 (n511, N116, n409);
nand U400 (n530, N139, n404);
nand U401 (n529, N103, n406);
nand U402 (n532, N127, n407);
nand U403 (n531, N115, n409);
nand U404 (n534, N138, n404);
nand U405 (n533, N102, n406);
nand U406 (n536, N126, n407);
nand U407 (n535, N114, n409);
nor U408 (N3671, n733, N37);
nand U409 (n556, N89, n414);
nand U410 (n555, N76, n416);
nand U411 (n558, N51, n418);
nand U412 (n557, N63, n419);
nand U413 (n560, N90, n414);
nand U414 (n559, N77, n416);
nand U415 (n562, N52, n418);
nand U416 (n561, N64, n419);
nand U417 (n580, N93, n414);
nand U418 (n579, N80, n416);
nand U419 (n582, N55, n418);
nand U420 (n581, N67, n419);
nand U421 (n584, N81, n414);
nand U422 (n583, N68, n416);
nand U423 (n586, N43, n418);
nand U424 (n585, N56, n419);
nand U425 (n588, N91, n414);
nand U426 (n587, N78, n416);
nand U427 (n590, N53, n418);
nand U428 (n589, N65, n419);
nand U429 (n592, N92, n414);
nand U430 (n591, N79, n416);
nand U431 (n594, N54, n418);
nand U432 (n593, N66, n419);
nand U433 (n564, N85, n414);
nand U434 (n563, N72, n416);
nand U435 (n566, N47, n418);
nand U436 (n565, N60, n419);
nand U437 (n568, N86, n414);
nand U438 (n567, N73, n416);
nand U439 (n570, N48, n418);
nand U440 (n569, N61, n419);
nand U441 (n571, N49, n418);
nand U442 (n574, N87, n415);
nand U443 (n573, N74, N234);
nand U444 (n576, N88, n414);
nand U445 (n575, N75, n416);
nand U446 (n578, N50, n418);
nand U447 (n577, N62, n419);
nand U448 (n742, n740, n828);
nand U449 (n743, n737, n829);
not U450 (n830, n741);
nor U451 (N3809, n831, N37);
nand U452 (n754, n752, n832);
nand U453 (n755, n749, n833);
nand U454 (n725, n723, n834);
nand U455 (n726, n720, n835);
nand U456 (n656, N14, n836);
not U457 (N2925, n656);
nand U458 (n432, N325, n296);
nand U459 (n431, N231, n295);
not U460 (N1726, n430);
not U461 (n837, n349);
nand U462 (n838, n659, n837);
nand U463 (n667, n660, n837);
nand U464 (n668, n661, n837);
nand U465 (n839, n399, n436);
nand U466 (n361, n764, n839);
nand U467 (n360, n840, n336);
nand U468 (n366, n663, n841);
nand U469 (n365, n363, N1821);
not U470 (n396, n364);
nand U471 (n842, n670, n668);
nand U472 (n843, n308, n425);
nand U473 (n844, n843, n842);
nand U474 (n845, n844, n667);
nand U475 (n846, n455, n845);
nand U476 (n847, n669, n848);
nand U477 (n849, n837, n846);
nand U478 (n850, n849, n847);
nand U479 (n289, n658, n837);
nand U480 (n288, n850, n838);
not U481 (n851, n438);
nand U482 (n293, N1, N3);
not U483 (N1448, N1277);
not U484 (n297, N1028);
nand U485 (n852, n359, n284);
nand U486 (n665, n368, n369);
nand U487 (n841, n767, n852);
nand U488 (n664, n395, n396);
nand U489 (n397, n851, n441);
nand U490 (n609, N340, n853);
nand U491 (n608, N343, n854);
nor U492 (n612, n855, N337);
nand U493 (n856, N337, n855);
nand U494 (n857, n607, n610);
nor U495 (n614, n610, n607);
nand U496 (n858, N256, n715);
nand U497 (n859, N259, n714);
nand U498 (n835, n859, n858);
nand U499 (n860, N346, n717);
nand U500 (n861, N349, n716);
nand U501 (n834, n861, n860);
nand U502 (n618, N328, n862);
nand U503 (n617, N331, n863);
nor U504 (n864, n724, n616);
nand U505 (n620, n616, n724);
nor U506 (n865, n613, n619);
nand U507 (n866, n619, n613);
nand U508 (n836, n866, n867);
nor U509 (n551, n868, n314);
nor U510 (n550, n410, n311);
nand U511 (n539, n301, n412);
nand U512 (n538, N1816, n727);
nor U513 (n542, n728, n537);
nor U514 (n541, n869, N1817);
not U515 (n870, n540);
nand U516 (n545, n308, n729);
nand U517 (n544, n320, n413);
nor U518 (n548, n730, n543);
nor U519 (n547, n871, N1818);
nor U520 (n448, n540, n872);
nor U521 (n447, n546, n870);
nand U522 (n554, n446, n317);
nand U523 (n553, n873, n411);
nand U524 (n603, N2012, N1820);
nand U525 (n602, N2014, N1821);
nand U526 (n874, N2020, n281);
nand U527 (n875, N2022, n282);
nand U528 (n829, n875, n874);
nand U529 (n876, N2016, n283);
nand U530 (n877, N2018, N1819);
nand U531 (n828, n877, n876);
nand U532 (n597, n329, n421);
nand U533 (n596, n294, n420);
nand U534 (n600, n399, n284);
nand U535 (n599, n336, N2010);
nand U536 (n878, n595, n879);
nor U537 (n450, n879, n595);
nand U538 (n880, n830, n449);
nor U539 (n605, n449, n830);
nand U540 (n881, n601, n604);
nor U541 (n882, n604, n601);
nor U542 (n831, n882, n883);
nand U543 (n639, N313, n291);
nand U544 (n638, N316, n744);
nand U545 (n642, N305, n402);
nand U546 (n641, N309, n403);
nand U547 (n645, n637, n884);
nand U548 (n644, n640, n885);
nand U549 (n648, N297, n400);
nand U550 (n647, N301, n401);
nor U551 (n651, n422, N355);
nor U552 (n650, n886, N294);
nand U553 (n887, n646, n649);
nor U554 (n653, n649, n646);
nand U555 (n888, n643, n652);
nor U556 (n889, n652, n643);
nor U557 (N2970, n889, n890);
nand U558 (n624, N272, n423);
nand U559 (n623, N275, n745);
nand U560 (n627, N266, n746);
nand U561 (n626, N269, n424);
nor U562 (n630, n891, n625);
nand U563 (n892, n625, n891);
nand U564 (n893, N284, n426);
nand U565 (n894, N287, n425);
nand U566 (n833, n894, n893);
nand U567 (n895, N278, n428);
nand U568 (n896, N281, n427);
nand U569 (n832, n896, n895);
nand U570 (n633, N263, n897);
nand U571 (n632, N352, n429);
nor U572 (n898, n753, n631);
nand U573 (n635, n631, n753);
nor U574 (n899, n628, n634);
nand U575 (n452, n634, n628);
nand U576 (n488, N269, n434);
nand U577 (n487, n756, N305);
nand U578 (n486, n756, n400);
nand U579 (n485, n424, n434);
nand U580 (n673, n830, n851);
nand U581 (n672, n438, n741);
nor U582 (n900, n449, n671);
nand U583 (n901, n671, n449);
nand U584 (n902, n901, n903);
nand U585 (n490, n420, n768);
nand U586 (n489, N246, n902);
nand U587 (n676, n294, n399);
nand U588 (n675, n336, n421);
nand U589 (n904, n905, n438);
nand U590 (n906, n674, n851);
nand U591 (n770, n906, n904);
nand U592 (n493, N25, n774);
nand U593 (n492, N29, n413);
nand U594 (n907, n908, N284);
nand U595 (n909, n491, n425);
nand U596 (n711, n909, n907);
nand U597 (n456, N287, n410);
nand U598 (n455, n314, n426);
nand U599 (n459, N294, n411);
nand U600 (n458, n317, n422);
nand U601 (n462, N301, n730);
nand U602 (n461, N1818, n400);
nand U603 (n465, N305, n412);
nand U604 (n464, N1816, n403);
nand U605 (n468, N297, n729);
nand U606 (n467, n320, n401);
nand U607 (n910, N263, n911);
nand U608 (n912, N20, n429);
nand U609 (n692, n912, n910);
nand U610 (n913, N256, n914);
nand U611 (n915, N19, n714);
nand U612 (n691, n915, n913);
nand U613 (n471, N256, n421);
nand U614 (n470, n294, n714);
nand U615 (n474, N269, N2014);
nand U616 (n473, n746, N1820);
nand U617 (n477, N266, N2012);
nand U618 (n476, n424, N1821);
nand U619 (n355, N275, N2018);
nand U620 (n375, n423, n283);
nand U621 (n481, N272, N2016);
nand U622 (n480, n745, N1819);
nand U623 (n350, N281, N2022);
nand U624 (n483, n428, n281);
nand U625 (n353, N278, N2020);
nand U626 (n379, n427, n282);
nand U627 (n495, n421, n768);
nand U628 (n494, N246, n851);
nand U629 (n497, N246, N2014);
nand U630 (n496, N2010, n768);
nand U631 (n499, N246, N2012);
nand U632 (n498, n399, n768);
not U633 (n300, n500);
not U634 (n408, N322);
not U635 (n848, n666);
not U636 (n440, N224);
not U637 (n867, n865);
not U638 (n621, n864);
not U639 (n890, n888);
not U640 (n615, n857);
not U641 (n654, n887);
not U642 (n883, n881);
not U643 (n734, n731);
not U644 (n453, n899);
not U645 (n636, n898);
not U646 (n891, n622);
not U647 (n885, n637);
not U648 (n863, N328);
not U649 (n855, N334);
not U650 (n854, N340);
not U651 (n879, n598);
not U652 (n903, n900);
not U653 (n897, N352);
not U654 (n629, n892);
not U655 (n886, N355);
not U656 (n884, n640);
not U657 (n862, N331);
not U658 (n611, n856);
not U659 (n853, N343);
not U660 (n417, N234);
not U661 (n451, n878);
not U662 (n606, n880);
not U663 (n871, n543);
not U664 (n869, n537);
not U665 (n872, n546);
not U666 (n873, n446);
not U667 (n868, n311);
not U668 (n757, n347);
not U669 (n840, n436);
not U670 (n905, n674);
not U671 (n772, n769);
not U672 (n908, n491);
not U673 (n802, N5);
not U674 (n805, N21);
not U675 (n799, N4);
not U676 (n914, N19);
not U677 (n911, N20);
not U678 (n814, N6);
not U679 (n817, N24);
not U680 (n808, N22);
not U681 (n811, N23);
not U682 (n783, N33);
not U683 (n786, N35);
not U684 (n777, N32);
not U685 (n780, N26);
not U686 (n789, N27);
not U687 (n792, N34);
endmodule