module c5315 (N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610, N613, N616, N619, N625, N631, N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128);
input N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610, N613, N616, N619, N625, N631;
output N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128;
wire N1042, N1043, N1067, N1080, N1092, N1104, N1146, N1148, N1149, N1150, N1151, N1156, N1157, N1161, N1173, N1185, N1197, N1209, N1213, N1216, N1219, N1223, N1235, N1247, N1259, N1271, N1280, N1292, N1303, N1315, N1327, N1339, N1351, N1363, N1375, N1378, N1381, N1384, N1387, N1390, N1393, N1396, N1415, N1418, N1421, N1424, N1427, N1430, N1433, N1436, N1455, N1462, N1469, N1475, N1479, N1482, N1492, N1495, N1498, N1501, N1504, N1507, N1510, N1513, N1516, N1519, N1522, N1525, N1542, N1545, N1548, N1551, N1554, N1557, N1560, N1563, N1566, N1573, N1580, N1583, N1588, N1594, N1597, N1600, N1603, N1606, N1609, N1612, N1615, N1618, N1621, N1624, N1627, N1630, N1633, N1636, N1639, N1642, N1645, N1648, N1651, N1654, N1657, N1660, N1663, N1675, N1685, N1697, N1709, N1721, N1727, N1731, N1743, N1755, N1758, N1761, N1769, N1777, N1785, N1793, N1800, N1807, N1814, N1821, N1824, N1827, N1830, N1833, N1836, N1839, N1842, N1845, N1848, N1851, N1854, N1857, N1860, N1863, N1866, N1869, N1872, N1875, N1878, N1881, N1884, N1887, N1890, N1893, N1896, N1899, N1902, N1905, N1908, N1911, N1914, N1917, N1920, N1923, N1926, N1929, N1932, N1935, N1938, N1941, N1944, N1947, N1950, N1953, N1956, N1959, N1962, N1965, N1968, N2349, N2350, N2585, N2586, N2587, N2588, N2589, N2591, N2592, N2593, N2594, N2595, N2596, N2597, N2598, N2599, N2600, N2601, N2602, N2603, N2604, N2605, N2606, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2614, N2615, N2616, N2617, N2618, N2619, N2620, N2621, N2622, N2624, N2625, N2626, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634, N2635, N2636, N2637, N2638, N2639, N2640, N2641, N2642, N2643, N2644, N2645, N2646, N2647, N2653, N2664, N2675, N2681, N2692, N2703, N2704, N2709, N2710, N2711, N2712, N2713, N2714, N2715, N2716, N2717, N2718, N2719, N2720, N2721, N2722, N2728, N2739, N2750, N2756, N2767, N2778, N2779, N2790, N2801, N2812, N2823, N2824, N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834, N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844, N2845, N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855, N2861, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875, N2876, N2877, N2882, N2891, N2901, N2902, N2903, N2904, N2905, N2906, N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2948, N2954, N2955, N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2969, N2970, N2971, N2972, N2973, N2974, N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3003, N3006, N3007, N3010, N3013, N3014, N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3038, N3041, N3052, N3063, N3068, N3071, N3072, N3073, N3074, N3075, N3086, N3097, N3108, N3119, N3130, N3141, N3142, N3143, N3144, N3145, N3146, N3147, N3158, N3169, N3180, N3191, N3194, N3195, N3196, N3197, N3198, N3199, N3200, N3203, N3401, N3402, N3403, N3404, N3405, N3406, N3407, N3408, N3409, N3410, N3411, N3412, N3413, N3414, N3415, N3416, N3444, N3445, N3446, N3447, N3448, N3449, N3450, N3451, N3452, N3453, N3454, N3455, N3456, N3459, N3460, N3461, N3462, N3463, N3464, N3465, N3466, N3481, N3482, N3483, N3484, N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509, N3510, N3511, N3512, N3513, N3514, N3515, N3558, N3559, N3560, N3561, N3562, N3563, N3605, N3606, N3607, N3608, N3609, N3610, N3614, N3615, N3616, N3617, N3618, N3619, N3620, N3621, N3622, N3623, N3624, N3625, N3626, N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3636, N3637, N3638, N3639, N3640, N3641, N3642, N3643, N3644, N3645, N3646, N3647, N3648, N3649, N3650, N3651, N3652, N3653, N3654, N3655, N3656, N3657, N3658, N3659, N3660, N3661, N3662, N3663, N3664, N3665, N3666, N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676, N3677, N3678, N3679, N3680, N3681, N3682, N3683, N3684, N3685, N3686, N3687, N3688, N3689, N3691, N3700, N3701, N3702, N3703, N3704, N3705, N3708, N3709, N3710, N3711, N3712, N3713, N3715, N3716, N3717, N3718, N3719, N3720, N3721, N3722, N3723, N3724, N3725, N3726, N3727, N3728, N3729, N3730, N3731, N3732, N3738, N3739, N3740, N3741, N3742, N3743, N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752, N3753, N3754, N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762, N3763, N3764, N3765, N3766, N3767, N3768, N3769, N3770, N3771, N3775, N3779, N3780, N3781, N3782, N3783, N3784, N3785, N3786, N3787, N3788, N3789, N3793, N3797, N3800, N3801, N3802, N3803, N3804, N3805, N3806, N3807, N3808, N3809, N3810, N3813, N3816, N3819, N3822, N3823, N3824, N3827, N3828, N3829, N3830, N3831, N3834, N3835, N3836, N3837, N3838, N3839, N3840, N3841, N3842, N3849, N3855, N3861, N3867, N3873, N3881, N3887, N3893, N3908, N3909, N3911, N3914, N3915, N3916, N3917, N3918, N3919, N3920, N3921, N3927, N3933, N3942, N3948, N3956, N3962, N3968, N3975, N3976, N3977, N3978, N3979, N3980, N3981, N3982, N3983, N3984, N3987, N3988, N3989, N3990, N3991, N3998, N4008, N4011, N4021, N4024, N4027, N4031, N4032, N4033, N4034, N4035, N4036, N4037, N4038, N4039, N4040, N4041, N4042, N4067, N4080, N4088, N4091, N4094, N4097, N4100, N4103, N4106, N4109, N4144, N4147, N4150, N4153, N4156, N4159, N4183, N4184, N4185, N4186, N4188, N4191, N4196, N4197, N4198, N4199, N4200, N4203, N4206, N4209, N4212, N4215, N4219, N4223, N4224, N4225, N4228, N4231, N4234, N4237, N4240, N4243, N4246, N4249, N4252, N4255, N4258, N4263, N4264, N4267, N4268, N4269, N4270, N4271, N4273, N4274, N4276, N4277, N4280, N4284, N4290, N4297, N4298, N4301, N4305, N4310, N4316, N4320, N4325, N4331, N4332, N4336, N4342, N4349, N4357, N4364, N4375, N4379, N4385, N4392, N4396, N4400, N4405, N4412, N4418, N4425, N4436, N4440, N4445, N4451, N4456, N4462, N4469, N4477, N4512, N4515, N4516, N4521, N4523, N4524, N4532, N4547, N4548, N4551, N4554, N4557, N4560, N4563, N4566, N4569, N4572, N4575, N4578, N4581, N4584, N4587, N4590, N4593, N4596, N4599, N4602, N4605, N4608, N4611, N4614, N4617, N4621, N4624, N4627, N4630, N4633, N4637, N4640, N4643, N4646, N4649, N4652, N4655, N4658, N4662, N4665, N4668, N4671, N4674, N4677, N4680, N4683, N4686, N4689, N4692, N4695, N4698, N4701, N4702, N4720, N4721, N4724, N4725, N4726, N4727, N4728, N4729, N4730, N4731, N4732, N4733, N4734, N4735, N4736, N4741, N4855, N4856, N4908, N4909, N4939, N4942, N4947, N4953, N4954, N4955, N4956, N4957, N4958, N4959, N4960, N4961, N4965, N4966, N4967, N4968, N4972, N4973, N4974, N4975, N4976, N4977, N4978, N4979, N4980, N4981, N4982, N4983, N4984, N4985, N4986, N4987, N5049, N5052, N5053, N5054, N5055, N5056, N5057, N5058, N5059, N5060, N5061, N5062, N5063, N5065, N5066, N5067, N5068, N5069, N5070, N5071, N5072, N5073, N5074, N5075, N5076, N5077, N5078, N5079, N5080, N5081, N5082, N5083, N5084, N5085, N5086, N5087, N5088, N5089, N5090, N5091, N5092, N5093, N5094, N5095, N5096, N5097, N5098, N5099, N5100, N5101, N5102, N5103, N5104, N5105, N5106, N5107, N5108, N5109, N5110, N5111, N5112, N5113, N5114, N5115, N5116, N5117, N5118, N5119, N5120, N5121, N5122, N5123, N5124, N5125, N5126, N5127, N5128, N5129, N5130, N5131, N5132, N5133, N5135, N5136, N5137, N5138, N5139, N5140, N5141, N5142, N5143, N5144, N5145, N5146, N5147, N5148, N5150, N5153, N5154, N5155, N5156, N5157, N5160, N5161, N5162, N5163, N5164, N5165, N5166, N5169, N5172, N5173, N5176, N5177, N5180, N5183, N5186, N5189, N5192, N5195, N5198, N5199, N5202, N5205, N5208, N5211, N5214, N5217, N5220, N5223, N5224, N5225, N5226, N5227, N5228, N5229, N5230, N5232, N5233, N5234, N5235, N5236, N5239, N5241, N5242, N5243, N5244, N5245, N5246, N5247, N5248, N5249, N5250, N5252, N5253, N5254, N5255, N5256, N5257, N5258, N5259, N5260, N5261, N5262, N5263, N5264, N5274, N5275, N5282, N5283, N5284, N5298, N5299, N5300, N5303, N5304, N5305, N5306, N5307, N5308, N5309, N5310, N5311, N5312, N5315, N5319, N5324, N5328, N5331, N5332, N5346, N5363, N5364, N5365, N5366, N5367, N5368, N5369, N5370, N5371, N5374, N5377, N5382, N5385, N5389, N5396, N5407, N5418, N5424, N5431, N5441, N5452, N5462, N5469, N5470, N5477, N5488, N5498, N5506, N5520, N5536, N5549, N5555, N5562, N5573, N5579, N5595, N5606, N5616, N5617, N5618, N5619, N5620, N5621, N5622, N5624, N5634, N5655, N5671, N5684, N5690, N5691, N5692, N5696, N5700, N5703, N5707, N5711, N5726, N5727, N5728, N5730, N5731, N5732, N5733, N5734, N5735, N5736, N5739, N5742, N5745, N5755, N5756, N5954, N5955, N5956, N6005, N6006, N6023, N6024, N6025, N6028, N6031, N6034, N6037, N6040, N6044, N6045, N6048, N6051, N6054, N6065, N6066, N6067, N6068, N6069, N6071, N6072, N6073, N6074, N6075, N6076, N6077, N6078, N6079, N6080, N6083, N6084, N6085, N6086, N6087, N6088, N6089, N6090, N6091, N6094, N6095, N6096, N6097, N6098, N6099, N6100, N6101, N6102, N6103, N6104, N6105, N6106, N6107, N6108, N6111, N6112, N6113, N6114, N6115, N6116, N6117, N6120, N6121, N6122, N6123, N6124, N6125, N6126, N6127, N6128, N6129, N6130, N6131, N6132, N6133, N6134, N6135, N6136, N6137, N6138, N6139, N6140, N6143, N6144, N6145, N6146, N6147, N6148, N6149, N6152, N6153, N6154, N6155, N6156, N6157, N6158, N6159, N6160, N6161, N6162, N6163, N6164, N6168, N6171, N6172, N6173, N6174, N6175, N6178, N6179, N6180, N6181, N6182, N6183, N6184, N6185, N6186, N6187, N6188, N6189, N6190, N6191, N6192, N6193, N6194, N6197, N6200, N6203, N6206, N6209, N6212, N6215, N6218, N6221, N6234, N6235, N6238, N6241, N6244, N6247, N6250, N6253, N6256, N6259, N6262, N6265, N6268, N6271, N6274, N6277, N6280, N6283, N6286, N6289, N6292, N6295, N6298, N6301, N6304, N6307, N6310, N6313, N6316, N6319, N6322, N6325, N6328, N6331, N6335, N6338, N6341, N6344, N6347, N6350, N6353, N6356, N6359, N6364, N6367, N6370, N6373, N6374, N6375, N6376, N6377, N6378, N6382, N6386, N6388, N6392, N6397, N6411, N6415, N6419, N6427, N6434, N6437, N6441, N6445, N6448, N6449, N6466, N6469, N6470, N6471, N6472, N6473, N6474, N6475, N6476, N6477, N6478, N6482, N6486, N6490, N6494, N6500, N6504, N6508, N6512, N6516, N6526, N6536, N6539, N6553, N6556, N6566, N6569, N6572, N6575, N6580, N6584, N6587, N6592, N6599, N6606, N6609, N6619, N6622, N6630, N6631, N6632, N6633, N6634, N6637, N6640, N6650, N6651, N6653, N6655, N6657, N6659, N6660, N6661, N6662, N6663, N6664, N6666, N6668, N6670, N6672, N6675, N6680, N6681, N6682, N6683, N6689, N6690, N6691, N6692, N6693, N6695, N6698, N6699, N6700, N6703, N6708, N6709, N6710, N6711, N6712, N6713, N6714, N6715, N6718, N6719, N6720, N6721, N6722, N6724, N6739, N6740, N6741, N6744, N6745, N6746, N6751, N6752, N6753, N6754, N6755, N6760, N6761, N6762, N6772, N6773, N6776, N6777, N6782, N6783, N6784, N6785, N6790, N6791, N6792, N6795, N6801, N6802, N6803, N6804, N6805, N6806, N6807, N6808, N6809, N6810, N6811, N6812, N6813, N6814, N6815, N6816, N6817, N6823, N6824, N6825, N6826, N6827, N6828, N6829, N6830, N6831, N6834, N6835, N6836, N6837, N6838, N6839, N6840, N6841, N6842, N6843, N6844, N6850, N6851, N6852, N6853, N6854, N6855, N6856, N6857, N6860, N6861, N6862, N6863, N6866, N6872, N6873, N6874, N6875, N6876, N6879, N6880, N6881, N6884, N6885, N6888, N6889, N6890, N6891, N6894, N6895, N6896, N6897, N6900, N6901, N6904, N6905, N6908, N6909, N6912, N6913, N6914, N6915, N6916, N6919, N6922, N6923, N6930, N6932, N6935, N6936, N6937, N6938, N6939, N6940, N6946, N6947, N6948, N6949, N6953, N6954, N6955, N6956, N6957, N6958, N6964, N6965, N6966, N6967, N6973, N6974, N6975, N6976, N6977, N6978, N6979, N6987, N6990, N6999, N7002, N7003, N7006, N7011, N7012, N7013, N7016, N7018, N7019, N7020, N7021, N7022, N7023, N7028, N7031, N7034, N7037, N7040, N7041, N7044, N7045, N7046, N7047, N7048, N7049, N7054, N7057, N7060, N7064, N7065, N7072, N7073, N7074, N7075, N7076, N7079, N7080, N7083, N7084, N7085, N7086, N7087, N7088, N7089, N7090, N7093, N7094, N7097, N7101, N7105, N7110, N7114, N7115, N7116, N7125, N7126, N7127, N7130, N7131, N7139, N7140, N7141, N7146, N7147, N7149, N7150, N7151, N7152, N7153, N7158, N7159, N7160, N7166, N7167, N7168, N7169, N7170, N7171, N7172, N7173, N7174, N7175, N7176, N7177, N7178, N7179, N7180, N7181, N7182, N7183, N7184, N7185, N7186, N7187, N7188, N7189, N7190, N7196, N7197, N7198, N7204, N7205, N7206, N7207, N7208, N7209, N7212, N7215, N7216, N7217, N7218, N7219, N7222, N7225, N7228, N7229, N7236, N7239, N7242, N7245, N7250, N7257, N7260, N7263, N7268, N7269, N7270, N7276, N7282, N7288, N7294, N7300, N7301, N7304, N7310, N7320, N7321, N7328, N7338, N7339, N7340, N7341, N7342, N7349, N7357, N7364, N7394, N7397, N7402, N7405, N7406, N7407, N7408, N7409, N7412, N7415, N7416, N7417, N7418, N7419, N7420, N7421, N7424, N7425, N7426, N7427, N7428, N7429, N7430, N7431, N7433, N7434, N7435, N7436, N7437, N7438, N7439, N7440, N7441, N7442, N7443, N7444, N7445, N7446, N7447, N7448, N7450, N7451, N7452, N7453, N7454, N7455, N7456, N7457, N7458, N7459, N7460, N7461, N7462, N7463, N7464, N7468, N7479, N7481, N7482, N7483, N7484, N7485, N7486, N7487, N7488, N7489, N7492, N7493, N7498, N7499, N7500, N7505, N7507, N7508, N7509, N7510, N7512, N7513, N7514, N7525, N7526, N7527, N7528, N7529, N7530, N7531, N7537, N7543, N7549, N7555, N7561, N7567, N7573, N7579, N7582, N7585, N7586, N7587, N7588, N7589, N7592, N7595, N7598, N7599, N7624, N7625, N7631, N7636, N7657, N7658, N7665, N7666, N7667, N7668, N7669, N7670, N7671, N7672, N7673, N7674, N7675, N7676, N7677, N7678, N7679, N7680, N7681, N7682, N7683, N7684, N7685, N7686, N7687, N7688, N7689, N7690, N7691, N7692, N7693, N7694, N7695, N7696, N7697, N7708, N7709, N7710, N7711, N7712, N7715, N7718, N7719, N7720, N7721, N7722, N7723, N7724, N7727, N7728, N7729, N7730, N7731, N7732, N7733, N7734, N7743, N7744, N7749, N7750, N7751, N7762, N7765, N7768, N7769, N7770, N7771, N7772, N7775, N7778, N7781, N7782, N7787, N7788, N7795, N7796, N7797, N7798, N7799, N7800, N7803, N7806, N7807, N7808, N7809, N7810, N7811, N7812, N7815, N7816, N7821, N7822, N7823, N7826, N7829, N7832, N7833, N7834, N7835, N7836, N7839, N7842, N7845, N7846, N7851, N7852, N7859, N7860, N7861, N7862, N7863, N7864, N7867, N7870, N7871, N7872, N7873, N7874, N7875, N7876, N7879, N7880, N7885, N7886, N7887, N7890, N7893, N7896, N7897, N7898, N7899, N7900, N7903, N7906, N7909, N7910, N7917, N7918, N7923, N7924, N7925, N7926, N7927, N7928, N7929, N7930, N7931, N7932, N7935, N7938, N7939, N7940, N7943, N7944, N7945, N7946, N7951, N7954, N7957, N7960, N7963, N7966, N7967, N7968, N7969, N7970, N7973, N7974, N7984, N7985, N7987, N7988, N7989, N7990, N7991, N7992, N7993, N7994, N7995, N7996, N7997, N7998, N8001, N8004, N8009, N8013, N8017, N8020, N8021, N8022, N8023, N8025, N8026, N8027, N8031, N8032, N8033, N8034, N8035, N8036, N8037, N8038, N8039, N8040, N8041, N8042, N8043, N8044, N8045, N8048, N8055, N8056, N8057, N8058, N8059, N8060, N8061, N8064, N8071, N8072, N8073, N8074, N8077, N8078, N8079, N8082, N8089, N8090, N8091, N8092, N8093, N8096, N8099, N8102, N8113, N8114, N8115, N8116, N8117, N8118, N8119, N8120, N8121, N8122, N8125, N8126;

buff U1 (N709,N141);
buff U2 (N816,N293);
and U3 (N1042,N135,N631);
not U4 (N1043,N591);
buff U5 (N1066,N592);
not U6 (N1067,N595);
not U7 (N1080,N596);
not U8 (N1092,N597);
not U9 (N1104,N598);
not U10 (N1137,N545);
not U11 (N1138,N348);
not U12 (N1139,N366);
and U13 (N1140,N552,N562);
not U14 (N1141,N549);
not U15 (N1142,N545);
not U16 (N1143,N545);
not U17 (N1144,N338);
not U18 (N1145,N358);
nand U19 (N1146,N373,N1);
and U20 (N1147,N141,N145);
not U21 (N1148,N592);
not U22 (N1149,N1042);
and U23 (N1150,N1043,N27);
and U24 (N1151,N386,N556);
not U25 (N1152,N245);
not U26 (N1153,N552);
not U27 (N1154,N562);
not U28 (N1155,N559);
and U29 (N1156,N386,N559,N556,N552);
not U30 (N1157,N566);
buff U31 (N1161,N571);
buff U32 (N1173,N574);
buff U33 (N1185,N571);
buff U34 (N1197,N574);
buff U35 (N1209,N137);
buff U36 (N1213,N137);
buff U37 (N1216,N141);
not U38 (N1219,N583);
buff U39 (N1223,N577);
buff U40 (N1235,N580);
buff U41 (N1247,N577);
buff U42 (N1259,N580);
buff U43 (N1271,N254);
buff U44 (N1280,N251);
buff U45 (N1292,N251);
buff U46 (N1303,N248);
buff U47 (N1315,N248);
buff U48 (N1327,N610);
buff U49 (N1339,N607);
buff U50 (N1351,N613);
buff U51 (N1363,N616);
buff U52 (N1375,N210);
buff U53 (N1378,N210);
buff U54 (N1381,N218);
buff U55 (N1384,N218);
buff U56 (N1387,N226);
buff U57 (N1390,N226);
buff U58 (N1393,N234);
buff U59 (N1396,N234);
buff U60 (N1415,N257);
buff U61 (N1418,N257);
buff U62 (N1421,N265);
buff U63 (N1424,N265);
buff U64 (N1427,N273);
buff U65 (N1430,N273);
buff U66 (N1433,N281);
buff U67 (N1436,N281);
buff U68 (N1455,N335);
buff U69 (N1462,N335);
buff U70 (N1469,N206);
and U71 (N1475,N27,N31);
buff U72 (N1479,N1);
buff U73 (N1482,N588);
buff U74 (N1492,N293);
buff U75 (N1495,N302);
buff U76 (N1498,N308);
buff U77 (N1501,N308);
buff U78 (N1504,N316);
buff U79 (N1507,N316);
buff U80 (N1510,N324);
buff U81 (N1513,N324);
buff U82 (N1516,N341);
buff U83 (N1519,N341);
buff U84 (N1522,N351);
buff U85 (N1525,N351);
buff U86 (N1542,N257);
buff U87 (N1545,N257);
buff U88 (N1548,N265);
buff U89 (N1551,N265);
buff U90 (N1554,N273);
buff U91 (N1557,N273);
buff U92 (N1560,N281);
buff U93 (N1563,N281);
buff U94 (N1566,N332);
buff U95 (N1573,N332);
buff U96 (N1580,N549);
and U97 (N1583,N31,N27);
not U98 (N1588,N588);
buff U99 (N1594,N324);
buff U100 (N1597,N324);
buff U101 (N1600,N341);
buff U102 (N1603,N341);
buff U103 (N1606,N351);
buff U104 (N1609,N351);
buff U105 (N1612,N293);
buff U106 (N1615,N302);
buff U107 (N1618,N308);
buff U108 (N1621,N308);
buff U109 (N1624,N316);
buff U110 (N1627,N316);
buff U111 (N1630,N361);
buff U112 (N1633,N361);
buff U113 (N1636,N210);
buff U114 (N1639,N210);
buff U115 (N1642,N218);
buff U116 (N1645,N218);
buff U117 (N1648,N226);
buff U118 (N1651,N226);
buff U119 (N1654,N234);
buff U120 (N1657,N234);
not U121 (N1660,N324);
buff U122 (N1663,N242);
buff U123 (N1675,N242);
buff U124 (N1685,N254);
buff U125 (N1697,N610);
buff U126 (N1709,N607);
buff U127 (N1721,N625);
buff U128 (N1727,N619);
buff U129 (N1731,N613);
buff U130 (N1743,N616);
not U131 (N1755,N599);
not U132 (N1758,N603);
buff U133 (N1761,N619);
buff U134 (N1769,N625);
buff U135 (N1777,N619);
buff U136 (N1785,N625);
buff U137 (N1793,N619);
buff U138 (N1800,N625);
buff U139 (N1807,N619);
buff U140 (N1814,N625);
buff U141 (N1821,N299);
buff U142 (N1824,N446);
buff U143 (N1827,N457);
buff U144 (N1830,N468);
buff U145 (N1833,N422);
buff U146 (N1836,N435);
buff U147 (N1839,N389);
buff U148 (N1842,N400);
buff U149 (N1845,N411);
buff U150 (N1848,N374);
buff U151 (N1851,N4);
buff U152 (N1854,N446);
buff U153 (N1857,N457);
buff U154 (N1860,N468);
buff U155 (N1863,N435);
buff U156 (N1866,N389);
buff U157 (N1869,N400);
buff U158 (N1872,N411);
buff U159 (N1875,N422);
buff U160 (N1878,N374);
buff U161 (N1881,N479);
buff U162 (N1884,N490);
buff U163 (N1887,N503);
buff U164 (N1890,N514);
buff U165 (N1893,N523);
buff U166 (N1896,N534);
buff U167 (N1899,N54);
buff U168 (N1902,N479);
buff U169 (N1905,N503);
buff U170 (N1908,N514);
buff U171 (N1911,N523);
buff U172 (N1914,N534);
buff U173 (N1917,N490);
buff U174 (N1920,N361);
buff U175 (N1923,N369);
buff U176 (N1926,N341);
buff U177 (N1929,N351);
buff U178 (N1932,N308);
buff U179 (N1935,N316);
buff U180 (N1938,N293);
buff U181 (N1941,N302);
buff U182 (N1944,N281);
buff U183 (N1947,N289);
buff U184 (N1950,N265);
buff U185 (N1953,N273);
buff U186 (N1956,N234);
buff U187 (N1959,N257);
buff U188 (N1962,N218);
buff U189 (N1965,N226);
buff U190 (N1968,N210);
not U191 (N1972,N1146);
and U192 (N2054,N136,N1148);
not U193 (N2060,N1150);
not U194 (N2061,N1151);
buff U195 (N2139,N1209);
buff U196 (N2142,N1216);
buff U197 (N2309,N1479);
and U198 (N2349,N1104,N514);
or U199 (N2350,N1067,N514);
buff U200 (N2387,N1580);
buff U201 (N2527,N1821);
not U202 (N2584,N1580);
and U203 (N2585,N170,N1161,N1173);
and U204 (N2586,N173,N1161,N1173);
and U205 (N2587,N167,N1161,N1173);
and U206 (N2588,N164,N1161,N1173);
and U207 (N2589,N161,N1161,N1173);
nand U208 (N2590,N1475,N140);
and U209 (N2591,N185,N1185,N1197);
and U210 (N2592,N158,N1185,N1197);
and U211 (N2593,N152,N1185,N1197);
and U212 (N2594,N146,N1185,N1197);
and U213 (N2595,N170,N1223,N1235);
and U214 (N2596,N173,N1223,N1235);
and U215 (N2597,N167,N1223,N1235);
and U216 (N2598,N164,N1223,N1235);
and U217 (N2599,N161,N1223,N1235);
and U218 (N2600,N185,N1247,N1259);
and U219 (N2601,N158,N1247,N1259);
and U220 (N2602,N152,N1247,N1259);
and U221 (N2603,N146,N1247,N1259);
and U222 (N2604,N106,N1731,N1743);
and U223 (N2605,N61,N1327,N1339);
and U224 (N2606,N106,N1697,N1709);
and U225 (N2607,N49,N1697,N1709);
and U226 (N2608,N103,N1697,N1709);
and U227 (N2609,N40,N1697,N1709);
and U228 (N2610,N37,N1697,N1709);
and U229 (N2611,N20,N1327,N1339);
and U230 (N2612,N17,N1327,N1339);
and U231 (N2613,N70,N1327,N1339);
and U232 (N2614,N64,N1327,N1339);
and U233 (N2615,N49,N1731,N1743);
and U234 (N2616,N103,N1731,N1743);
and U235 (N2617,N40,N1731,N1743);
and U236 (N2618,N37,N1731,N1743);
and U237 (N2619,N20,N1351,N1363);
and U238 (N2620,N17,N1351,N1363);
and U239 (N2621,N70,N1351,N1363);
and U240 (N2622,N64,N1351,N1363);
not U241 (N2623,N1475);
and U242 (N2624,N123,N1758,N599);
and U243 (N2625,N1777,N1785);
and U244 (N2626,N61,N1351,N1363);
and U245 (N2627,N1761,N1769);
not U246 (N2628,N1824);
not U247 (N2629,N1827);
not U248 (N2630,N1830);
not U249 (N2631,N1833);
not U250 (N2632,N1836);
not U251 (N2633,N1839);
not U252 (N2634,N1842);
not U253 (N2635,N1845);
not U254 (N2636,N1848);
not U255 (N2637,N1851);
not U256 (N2638,N1854);
not U257 (N2639,N1857);
not U258 (N2640,N1860);
not U259 (N2641,N1863);
not U260 (N2642,N1866);
not U261 (N2643,N1869);
not U262 (N2644,N1872);
not U263 (N2645,N1875);
not U264 (N2646,N1878);
buff U265 (N2647,N1209);
not U266 (N2653,N1161);
not U267 (N2664,N1173);
buff U268 (N2675,N1209);
not U269 (N2681,N1185);
not U270 (N2692,N1197);
and U271 (N2703,N179,N1185,N1197);
buff U272 (N2704,N1479);
not U273 (N2709,N1881);
not U274 (N2710,N1884);
not U275 (N2711,N1887);
not U276 (N2712,N1890);
not U277 (N2713,N1893);
not U278 (N2714,N1896);
not U279 (N2715,N1899);
not U280 (N2716,N1902);
not U281 (N2717,N1905);
not U282 (N2718,N1908);
not U283 (N2719,N1911);
not U284 (N2720,N1914);
not U285 (N2721,N1917);
buff U286 (N2722,N1213);
not U287 (N2728,N1223);
not U288 (N2739,N1235);
buff U289 (N2750,N1213);
not U290 (N2756,N1247);
not U291 (N2767,N1259);
and U292 (N2778,N179,N1247,N1259);
not U293 (N2779,N1327);
not U294 (N2790,N1339);
not U295 (N2801,N1351);
not U296 (N2812,N1363);
not U297 (N2823,N1375);
not U298 (N2824,N1378);
not U299 (N2825,N1381);
not U300 (N2826,N1384);
not U301 (N2827,N1387);
not U302 (N2828,N1390);
not U303 (N2829,N1393);
not U304 (N2830,N1396);
and U305 (N2831,N1104,N457,N1378);
and U306 (N2832,N1104,N468,N1384);
and U307 (N2833,N1104,N422,N1390);
and U308 (N2834,N1104,N435,N1396);
and U309 (N2835,N1067,N1375);
and U310 (N2836,N1067,N1381);
and U311 (N2837,N1067,N1387);
and U312 (N2838,N1067,N1393);
not U313 (N2839,N1415);
not U314 (N2840,N1418);
not U315 (N2841,N1421);
not U316 (N2842,N1424);
not U317 (N2843,N1427);
not U318 (N2844,N1430);
not U319 (N2845,N1433);
not U320 (N2846,N1436);
and U321 (N2847,N1104,N389,N1418);
and U322 (N2848,N1104,N400,N1424);
and U323 (N2849,N1104,N411,N1430);
and U324 (N2850,N1104,N374,N1436);
and U325 (N2851,N1067,N1415);
and U326 (N2852,N1067,N1421);
and U327 (N2853,N1067,N1427);
and U328 (N2854,N1067,N1433);
not U329 (N2855,N1455);
not U330 (N2861,N1462);
and U331 (N2867,N292,N1455);
and U332 (N2868,N288,N1455);
and U333 (N2869,N280,N1455);
and U334 (N2870,N272,N1455);
and U335 (N2871,N264,N1455);
and U336 (N2872,N241,N1462);
and U337 (N2873,N233,N1462);
and U338 (N2874,N225,N1462);
and U339 (N2875,N217,N1462);
and U340 (N2876,N209,N1462);
buff U341 (N2877,N1216);
not U342 (N2882,N1482);
not U343 (N2891,N1475);
not U344 (N2901,N1492);
not U345 (N2902,N1495);
not U346 (N2903,N1498);
not U347 (N2904,N1501);
not U348 (N2905,N1504);
not U349 (N2906,N1507);
and U350 (N2907,N1303,N1495);
and U351 (N2908,N1303,N479,N1501);
and U352 (N2909,N1303,N490,N1507);
and U353 (N2910,N1663,N1492);
and U354 (N2911,N1663,N1498);
and U355 (N2912,N1663,N1504);
not U356 (N2913,N1510);
not U357 (N2914,N1513);
not U358 (N2915,N1516);
not U359 (N2916,N1519);
not U360 (N2917,N1522);
not U361 (N2918,N1525);
and U362 (N2919,N1104,N503,N1513);
not U363 (N2920,N2349);
and U364 (N2921,N1104,N523,N1519);
and U365 (N2922,N1104,N534,N1525);
and U366 (N2923,N1067,N1510);
and U367 (N2924,N1067,N1516);
and U368 (N2925,N1067,N1522);
not U369 (N2926,N1542);
not U370 (N2927,N1545);
not U371 (N2928,N1548);
not U372 (N2929,N1551);
not U373 (N2930,N1554);
not U374 (N2931,N1557);
not U375 (N2932,N1560);
not U376 (N2933,N1563);
and U377 (N2934,N1303,N389,N1545);
and U378 (N2935,N1303,N400,N1551);
and U379 (N2936,N1303,N411,N1557);
and U380 (N2937,N1303,N374,N1563);
and U381 (N2938,N1663,N1542);
and U382 (N2939,N1663,N1548);
and U383 (N2940,N1663,N1554);
and U384 (N2941,N1663,N1560);
not U385 (N2942,N1566);
not U386 (N2948,N1573);
and U387 (N2954,N372,N1566);
and U388 (N2955,N366,N1566);
and U389 (N2956,N358,N1566);
and U390 (N2957,N348,N1566);
and U391 (N2958,N338,N1566);
and U392 (N2959,N331,N1573);
and U393 (N2960,N323,N1573);
and U394 (N2961,N315,N1573);
and U395 (N2962,N307,N1573);
and U396 (N2963,N299,N1573);
not U397 (N2964,N1588);
and U398 (N2969,N83,N1588);
and U399 (N2970,N86,N1588);
and U400 (N2971,N88,N1588);
and U401 (N2972,N88,N1588);
not U402 (N2973,N1594);
not U403 (N2974,N1597);
not U404 (N2975,N1600);
not U405 (N2976,N1603);
not U406 (N2977,N1606);
not U407 (N2978,N1609);
and U408 (N2979,N1315,N503,N1597);
and U409 (N2980,N1315,N514);
and U410 (N2981,N1315,N523,N1603);
and U411 (N2982,N1315,N534,N1609);
and U412 (N2983,N1675,N1594);
or U413 (N2984,N1675,N514);
and U414 (N2985,N1675,N1600);
and U415 (N2986,N1675,N1606);
not U416 (N2987,N1612);
not U417 (N2988,N1615);
not U418 (N2989,N1618);
not U419 (N2990,N1621);
not U420 (N2991,N1624);
not U421 (N2992,N1627);
and U422 (N2993,N1315,N1615);
and U423 (N2994,N1315,N479,N1621);
and U424 (N2995,N1315,N490,N1627);
and U425 (N2996,N1675,N1612);
and U426 (N2997,N1675,N1618);
and U427 (N2998,N1675,N1624);
not U428 (N2999,N1630);
buff U429 (N3000,N1469);
buff U430 (N3003,N1469);
not U431 (N3006,N1633);
buff U432 (N3007,N1469);
buff U433 (N3010,N1469);
and U434 (N3013,N1315,N1630);
and U435 (N3014,N1315,N1633);
not U436 (N3015,N1636);
not U437 (N3016,N1639);
not U438 (N3017,N1642);
not U439 (N3018,N1645);
not U440 (N3019,N1648);
not U441 (N3020,N1651);
not U442 (N3021,N1654);
not U443 (N3022,N1657);
and U444 (N3023,N1303,N457,N1639);
and U445 (N3024,N1303,N468,N1645);
and U446 (N3025,N1303,N422,N1651);
and U447 (N3026,N1303,N435,N1657);
and U448 (N3027,N1663,N1636);
and U449 (N3028,N1663,N1642);
and U450 (N3029,N1663,N1648);
and U451 (N3030,N1663,N1654);
not U452 (N3031,N1920);
not U453 (N3032,N1923);
not U454 (N3033,N1926);
not U455 (N3034,N1929);
buff U456 (N3035,N1660);
buff U457 (N3038,N1660);
not U458 (N3041,N1697);
not U459 (N3052,N1709);
not U460 (N3063,N1721);
not U461 (N3068,N1727);
and U462 (N3071,N97,N1721);
and U463 (N3072,N94,N1721);
and U464 (N3073,N97,N1721);
and U465 (N3074,N94,N1721);
not U466 (N3075,N1731);
not U467 (N3086,N1743);
not U468 (N3097,N1761);
not U469 (N3108,N1769);
not U470 (N3119,N1777);
not U471 (N3130,N1785);
not U472 (N3141,N1944);
not U473 (N3142,N1947);
not U474 (N3143,N1950);
not U475 (N3144,N1953);
not U476 (N3145,N1956);
not U477 (N3146,N1959);
not U478 (N3147,N1793);
not U479 (N3158,N1800);
not U480 (N3169,N1807);
not U481 (N3180,N1814);
buff U482 (N3191,N1821);
not U483 (N3194,N1932);
not U484 (N3195,N1935);
not U485 (N3196,N1938);
not U486 (N3197,N1941);
not U487 (N3198,N1962);
not U488 (N3199,N1965);
buff U489 (N3200,N1469);
not U490 (N3203,N1968);
buff U491 (N3357,N2704);
buff U492 (N3358,N2704);
buff U493 (N3359,N2704);
buff U494 (N3360,N2704);
and U495 (N3401,N457,N1092,N2824);
and U496 (N3402,N468,N1092,N2826);
and U497 (N3403,N422,N1092,N2828);
and U498 (N3404,N435,N1092,N2830);
and U499 (N3405,N1080,N2823);
and U500 (N3406,N1080,N2825);
and U501 (N3407,N1080,N2827);
and U502 (N3408,N1080,N2829);
and U503 (N3409,N389,N1092,N2840);
and U504 (N3410,N400,N1092,N2842);
and U505 (N3411,N411,N1092,N2844);
and U506 (N3412,N374,N1092,N2846);
and U507 (N3413,N1080,N2839);
and U508 (N3414,N1080,N2841);
and U509 (N3415,N1080,N2843);
and U510 (N3416,N1080,N2845);
and U511 (N3444,N1280,N2902);
and U512 (N3445,N479,N1280,N2904);
and U513 (N3446,N490,N1280,N2906);
and U514 (N3447,N1685,N2901);
and U515 (N3448,N1685,N2903);
and U516 (N3449,N1685,N2905);
and U517 (N3450,N503,N1092,N2914);
and U518 (N3451,N523,N1092,N2916);
and U519 (N3452,N534,N1092,N2918);
and U520 (N3453,N1080,N2913);
and U521 (N3454,N1080,N2915);
and U522 (N3455,N1080,N2917);
and U523 (N3456,N2920,N2350);
and U524 (N3459,N389,N1280,N2927);
and U525 (N3460,N400,N1280,N2929);
and U526 (N3461,N411,N1280,N2931);
and U527 (N3462,N374,N1280,N2933);
and U528 (N3463,N1685,N2926);
and U529 (N3464,N1685,N2928);
and U530 (N3465,N1685,N2930);
and U531 (N3466,N1685,N2932);
and U532 (N3481,N503,N1292,N2974);
not U533 (N3482,N2980);
and U534 (N3483,N523,N1292,N2976);
and U535 (N3484,N534,N1292,N2978);
and U536 (N3485,N1271,N2973);
and U537 (N3486,N1271,N2975);
and U538 (N3487,N1271,N2977);
and U539 (N3488,N1292,N2988);
and U540 (N3489,N479,N1292,N2990);
and U541 (N3490,N490,N1292,N2992);
and U542 (N3491,N1271,N2987);
and U543 (N3492,N1271,N2989);
and U544 (N3493,N1271,N2991);
and U545 (N3502,N1292,N2999);
and U546 (N3503,N1292,N3006);
and U547 (N3504,N457,N1280,N3016);
and U548 (N3505,N468,N1280,N3018);
and U549 (N3506,N422,N1280,N3020);
and U550 (N3507,N435,N1280,N3022);
and U551 (N3508,N1685,N3015);
and U552 (N3509,N1685,N3017);
and U553 (N3510,N1685,N3019);
and U554 (N3511,N1685,N3021);
nand U555 (N3512,N1923,N3031);
nand U556 (N3513,N1920,N3032);
nand U557 (N3514,N1929,N3033);
nand U558 (N3515,N1926,N3034);
nand U559 (N3558,N1947,N3141);
nand U560 (N3559,N1944,N3142);
nand U561 (N3560,N1953,N3143);
nand U562 (N3561,N1950,N3144);
nand U563 (N3562,N1959,N3145);
nand U564 (N3563,N1956,N3146);
buff U565 (N3604,N3191);
nand U566 (N3605,N1935,N3194);
nand U567 (N3606,N1932,N3195);
nand U568 (N3607,N1941,N3196);
nand U569 (N3608,N1938,N3197);
nand U570 (N3609,N1965,N3198);
nand U571 (N3610,N1962,N3199);
not U572 (N3613,N3191);
and U573 (N3614,N2882,N2891);
and U574 (N3615,N1482,N2891);
and U575 (N3616,N200,N2653,N1173);
and U576 (N3617,N203,N2653,N1173);
and U577 (N3618,N197,N2653,N1173);
and U578 (N3619,N194,N2653,N1173);
and U579 (N3620,N191,N2653,N1173);
and U580 (N3621,N182,N2681,N1197);
and U581 (N3622,N188,N2681,N1197);
and U582 (N3623,N155,N2681,N1197);
and U583 (N3624,N149,N2681,N1197);
and U584 (N3625,N2882,N2891);
and U585 (N3626,N1482,N2891);
and U586 (N3627,N200,N2728,N1235);
and U587 (N3628,N203,N2728,N1235);
and U588 (N3629,N197,N2728,N1235);
and U589 (N3630,N194,N2728,N1235);
and U590 (N3631,N191,N2728,N1235);
and U591 (N3632,N182,N2756,N1259);
and U592 (N3633,N188,N2756,N1259);
and U593 (N3634,N155,N2756,N1259);
and U594 (N3635,N149,N2756,N1259);
and U595 (N3636,N2882,N2891);
and U596 (N3637,N1482,N2891);
and U597 (N3638,N109,N3075,N1743);
and U598 (N3639,N2882,N2891);
and U599 (N3640,N1482,N2891);
and U600 (N3641,N11,N2779,N1339);
and U601 (N3642,N109,N3041,N1709);
and U602 (N3643,N46,N3041,N1709);
and U603 (N3644,N100,N3041,N1709);
and U604 (N3645,N91,N3041,N1709);
and U605 (N3646,N43,N3041,N1709);
and U606 (N3647,N76,N2779,N1339);
and U607 (N3648,N73,N2779,N1339);
and U608 (N3649,N67,N2779,N1339);
and U609 (N3650,N14,N2779,N1339);
and U610 (N3651,N46,N3075,N1743);
and U611 (N3652,N100,N3075,N1743);
and U612 (N3653,N91,N3075,N1743);
and U613 (N3654,N43,N3075,N1743);
and U614 (N3655,N76,N2801,N1363);
and U615 (N3656,N73,N2801,N1363);
and U616 (N3657,N67,N2801,N1363);
and U617 (N3658,N14,N2801,N1363);
and U618 (N3659,N120,N3119,N1785);
and U619 (N3660,N11,N2801,N1363);
and U620 (N3661,N118,N3097,N1769);
and U621 (N3662,N176,N2681,N1197);
and U622 (N3663,N176,N2756,N1259);
or U623 (N3664,N2831,N3401);
or U624 (N3665,N2832,N3402);
or U625 (N3666,N2833,N3403);
or U626 (N3667,N2834,N3404);
or U627 (N3668,N2835,N3405,N457);
or U628 (N3669,N2836,N3406,N468);
or U629 (N3670,N2837,N3407,N422);
or U630 (N3671,N2838,N3408,N435);
or U631 (N3672,N2847,N3409);
or U632 (N3673,N2848,N3410);
or U633 (N3674,N2849,N3411);
or U634 (N3675,N2850,N3412);
or U635 (N3676,N2851,N3413,N389);
or U636 (N3677,N2852,N3414,N400);
or U637 (N3678,N2853,N3415,N411);
or U638 (N3679,N2854,N3416,N374);
and U639 (N3680,N289,N2855);
and U640 (N3681,N281,N2855);
and U641 (N3682,N273,N2855);
and U642 (N3683,N265,N2855);
and U643 (N3684,N257,N2855);
and U644 (N3685,N234,N2861);
and U645 (N3686,N226,N2861);
and U646 (N3687,N218,N2861);
and U647 (N3688,N210,N2861);
and U648 (N3689,N206,N2861);
not U649 (N3691,N2891);
or U650 (N3700,N2907,N3444);
or U651 (N3701,N2908,N3445);
or U652 (N3702,N2909,N3446);
or U653 (N3703,N2911,N3448,N479);
or U654 (N3704,N2912,N3449,N490);
or U655 (N3705,N2910,N3447);
or U656 (N3708,N2919,N3450);
or U657 (N3709,N2921,N3451);
or U658 (N3710,N2922,N3452);
or U659 (N3711,N2923,N3453,N503);
or U660 (N3712,N2924,N3454,N523);
or U661 (N3713,N2925,N3455,N534);
or U662 (N3715,N2934,N3459);
or U663 (N3716,N2935,N3460);
or U664 (N3717,N2936,N3461);
or U665 (N3718,N2937,N3462);
or U666 (N3719,N2938,N3463,N389);
or U667 (N3720,N2939,N3464,N400);
or U668 (N3721,N2940,N3465,N411);
or U669 (N3722,N2941,N3466,N374);
and U670 (N3723,N369,N2942);
and U671 (N3724,N361,N2942);
and U672 (N3725,N351,N2942);
and U673 (N3726,N341,N2942);
and U674 (N3727,N324,N2948);
and U675 (N3728,N316,N2948);
and U676 (N3729,N308,N2948);
and U677 (N3730,N302,N2948);
and U678 (N3731,N293,N2948);
or U679 (N3732,N2942,N2958);
and U680 (N3738,N83,N2964);
and U681 (N3739,N87,N2964);
and U682 (N3740,N34,N2964);
and U683 (N3741,N34,N2964);
or U684 (N3742,N2979,N3481);
or U685 (N3743,N2981,N3483);
or U686 (N3744,N2982,N3484);
or U687 (N3745,N2983,N3485,N503);
or U688 (N3746,N2985,N3486,N523);
or U689 (N3747,N2986,N3487,N534);
or U690 (N3748,N2993,N3488);
or U691 (N3749,N2994,N3489);
or U692 (N3750,N2995,N3490);
or U693 (N3751,N2997,N3492,N479);
or U694 (N3752,N2998,N3493,N490);
not U695 (N3753,N3000);
not U696 (N3754,N3003);
not U697 (N3755,N3007);
not U698 (N3756,N3010);
or U699 (N3757,N3013,N3502);
and U700 (N3758,N1315,N446,N3003);
or U701 (N3759,N3014,N3503);
and U702 (N3760,N1315,N446,N3010);
and U703 (N3761,N1675,N3000);
and U704 (N3762,N1675,N3007);
or U705 (N3763,N3023,N3504);
or U706 (N3764,N3024,N3505);
or U707 (N3765,N3025,N3506);
or U708 (N3766,N3026,N3507);
or U709 (N3767,N3027,N3508,N457);
or U710 (N3768,N3028,N3509,N468);
or U711 (N3769,N3029,N3510,N422);
or U712 (N3770,N3030,N3511,N435);
nand U713 (N3771,N3512,N3513);
nand U714 (N3775,N3514,N3515);
not U715 (N3779,N3035);
not U716 (N3780,N3038);
and U717 (N3781,N117,N3097,N1769);
and U718 (N3782,N126,N3097,N1769);
and U719 (N3783,N127,N3097,N1769);
and U720 (N3784,N128,N3097,N1769);
and U721 (N3785,N131,N3119,N1785);
and U722 (N3786,N129,N3119,N1785);
and U723 (N3787,N119,N3119,N1785);
and U724 (N3788,N130,N3119,N1785);
nand U725 (N3789,N3558,N3559);
nand U726 (N3793,N3560,N3561);
nand U727 (N3797,N3562,N3563);
and U728 (N3800,N122,N3147,N1800);
and U729 (N3801,N113,N3147,N1800);
and U730 (N3802,N53,N3147,N1800);
and U731 (N3803,N114,N3147,N1800);
and U732 (N3804,N115,N3147,N1800);
and U733 (N3805,N52,N3169,N1814);
and U734 (N3806,N112,N3169,N1814);
and U735 (N3807,N116,N3169,N1814);
and U736 (N3808,N121,N3169,N1814);
and U737 (N3809,N123,N3169,N1814);
nand U738 (N3810,N3607,N3608);
nand U739 (N3813,N3605,N3606);
and U740 (N3816,N3482,N2984);
or U741 (N3819,N2996,N3491);
not U742 (N3822,N3200);
nand U743 (N3823,N3200,N3203);
nand U744 (N3824,N3609,N3610);
not U745 (N3827,N3456);
or U746 (N3828,N3739,N2970);
or U747 (N3829,N3740,N2971);
or U748 (N3830,N3741,N2972);
or U749 (N3831,N3738,N2969);
not U750 (N3834,N3664);
not U751 (N3835,N3665);
not U752 (N3836,N3666);
not U753 (N3837,N3667);
not U754 (N3838,N3672);
not U755 (N3839,N3673);
not U756 (N3840,N3674);
not U757 (N3841,N3675);
or U758 (N3842,N3681,N2868);
or U759 (N3849,N3682,N2869);
or U760 (N3855,N3683,N2870);
or U761 (N3861,N3684,N2871);
or U762 (N3867,N3685,N2872);
or U763 (N3873,N3686,N2873);
or U764 (N3881,N3687,N2874);
or U765 (N3887,N3688,N2875);
or U766 (N3893,N3689,N2876);
not U767 (N3908,N3701);
not U768 (N3909,N3702);
not U769 (N3911,N3700);
not U770 (N3914,N3708);
not U771 (N3915,N3709);
not U772 (N3916,N3710);
not U773 (N3917,N3715);
not U774 (N3918,N3716);
not U775 (N3919,N3717);
not U776 (N3920,N3718);
or U777 (N3921,N3724,N2955);
or U778 (N3927,N3725,N2956);
or U779 (N3933,N3726,N2957);
or U780 (N3942,N3727,N2959);
or U781 (N3948,N3728,N2960);
or U782 (N3956,N3729,N2961);
or U783 (N3962,N3730,N2962);
or U784 (N3968,N3731,N2963);
not U785 (N3975,N3742);
not U786 (N3976,N3743);
not U787 (N3977,N3744);
not U788 (N3978,N3749);
not U789 (N3979,N3750);
and U790 (N3980,N446,N1292,N3754);
and U791 (N3981,N446,N1292,N3756);
and U792 (N3982,N1271,N3753);
and U793 (N3983,N1271,N3755);
not U794 (N3984,N3757);
not U795 (N3987,N3759);
not U796 (N3988,N3763);
not U797 (N3989,N3764);
not U798 (N3990,N3765);
not U799 (N3991,N3766);
and U800 (N3998,N3456,N3119,N3130);
or U801 (N4008,N3723,N2954);
or U802 (N4011,N3680,N2867);
not U803 (N4021,N3748);
nand U804 (N4024,N1968,N3822);
not U805 (N4027,N3705);
and U806 (N4031,N3828,N1583);
and U807 (N4032,N24,N2882,N3691);
and U808 (N4033,N25,N1482,N3691);
and U809 (N4034,N26,N2882,N3691);
and U810 (N4035,N81,N1482,N3691);
and U811 (N4036,N3829,N1583);
and U812 (N4037,N79,N2882,N3691);
and U813 (N4038,N23,N1482,N3691);
and U814 (N4039,N82,N2882,N3691);
and U815 (N4040,N80,N1482,N3691);
and U816 (N4041,N3830,N1583);
and U817 (N4042,N3831,N1583);
and U818 (N4067,N3732,N514);
and U819 (N4080,N514,N3732);
and U820 (N4088,N3834,N3668);
and U821 (N4091,N3835,N3669);
and U822 (N4094,N3836,N3670);
and U823 (N4097,N3837,N3671);
and U824 (N4100,N3838,N3676);
and U825 (N4103,N3839,N3677);
and U826 (N4106,N3840,N3678);
and U827 (N4109,N3841,N3679);
and U828 (N4144,N3908,N3703);
and U829 (N4147,N3909,N3704);
buff U830 (N4150,N3705);
and U831 (N4153,N3914,N3711);
and U832 (N4156,N3915,N3712);
and U833 (N4159,N3916,N3713);
or U834 (N4183,N3758,N3980);
or U835 (N4184,N3760,N3981);
or U836 (N4185,N3761,N3982,N446);
or U837 (N4186,N3762,N3983,N446);
not U838 (N4188,N3771);
not U839 (N4191,N3775);
and U840 (N4196,N3775,N3771,N3035);
and U841 (N4197,N3987,N3119,N3130);
and U842 (N4198,N3920,N3722);
not U843 (N4199,N3816);
not U844 (N4200,N3789);
not U845 (N4203,N3793);
buff U846 (N4206,N3797);
buff U847 (N4209,N3797);
buff U848 (N4212,N3732);
buff U849 (N4215,N3732);
buff U850 (N4219,N3732);
not U851 (N4223,N3810);
not U852 (N4224,N3813);
and U853 (N4225,N3918,N3720);
and U854 (N4228,N3919,N3721);
and U855 (N4231,N3991,N3770);
and U856 (N4234,N3917,N3719);
and U857 (N4237,N3989,N3768);
and U858 (N4240,N3990,N3769);
and U859 (N4243,N3988,N3767);
and U860 (N4246,N3976,N3746);
and U861 (N4249,N3977,N3747);
and U862 (N4252,N3975,N3745);
and U863 (N4255,N3978,N3751);
and U864 (N4258,N3979,N3752);
not U865 (N4263,N3819);
nand U866 (N4264,N4024,N3823);
not U867 (N4267,N3824);
and U868 (N4268,N446,N3893);
not U869 (N4269,N3911);
not U870 (N4270,N3984);
and U871 (N4271,N3893,N446);
not U872 (N4272,N4031);
or U873 (N4273,N4032,N4033,N3614,N3615);
or U874 (N4274,N4034,N4035,N3625,N3626);
not U875 (N4275,N4036);
or U876 (N4276,N4037,N4038,N3636,N3637);
or U877 (N4277,N4039,N4040,N3639,N3640);
not U878 (N4278,N4041);
not U879 (N4279,N4042);
and U880 (N4280,N3887,N457);
and U881 (N4284,N3881,N468);
and U882 (N4290,N422,N3873);
and U883 (N4297,N3867,N435);
and U884 (N4298,N3861,N389);
and U885 (N4301,N3855,N400);
and U886 (N4305,N3849,N411);
and U887 (N4310,N3842,N374);
and U888 (N4316,N457,N3887);
and U889 (N4320,N468,N3881);
and U890 (N4325,N422,N3873);
and U891 (N4331,N435,N3867);
and U892 (N4332,N389,N3861);
and U893 (N4336,N400,N3855);
and U894 (N4342,N411,N3849);
and U895 (N4349,N374,N3842);
not U896 (N4357,N3968);
not U897 (N4364,N3962);
buff U898 (N4375,N3962);
and U899 (N4379,N3956,N479);
and U900 (N4385,N490,N3948);
and U901 (N4392,N3942,N503);
and U902 (N4396,N3933,N523);
and U903 (N4400,N3927,N534);
not U904 (N4405,N3921);
buff U905 (N4412,N3921);
not U906 (N4418,N3968);
not U907 (N4425,N3962);
buff U908 (N4436,N3962);
and U909 (N4440,N479,N3956);
and U910 (N4445,N490,N3948);
and U911 (N4451,N503,N3942);
and U912 (N4456,N523,N3933);
and U913 (N4462,N534,N3927);
buff U914 (N4469,N3921);
not U915 (N4477,N3921);
buff U916 (N4512,N3968);
not U917 (N4515,N4183);
not U918 (N4516,N4184);
not U919 (N4521,N4008);
not U920 (N4523,N4011);
not U921 (N4524,N4198);
not U922 (N4532,N3984);
and U923 (N4547,N3911,N3169,N3180);
buff U924 (N4548,N3893);
buff U925 (N4551,N3887);
buff U926 (N4554,N3881);
buff U927 (N4557,N3873);
buff U928 (N4560,N3867);
buff U929 (N4563,N3861);
buff U930 (N4566,N3855);
buff U931 (N4569,N3849);
buff U932 (N4572,N3842);
nor U933 (N4575,N422,N3873);
buff U934 (N4578,N3893);
buff U935 (N4581,N3887);
buff U936 (N4584,N3881);
buff U937 (N4587,N3867);
buff U938 (N4590,N3861);
buff U939 (N4593,N3855);
buff U940 (N4596,N3849);
buff U941 (N4599,N3873);
buff U942 (N4602,N3842);
nor U943 (N4605,N422,N3873);
nor U944 (N4608,N374,N3842);
buff U945 (N4611,N3956);
buff U946 (N4614,N3948);
buff U947 (N4617,N3942);
buff U948 (N4621,N3933);
buff U949 (N4624,N3927);
nor U950 (N4627,N490,N3948);
buff U951 (N4630,N3956);
buff U952 (N4633,N3942);
buff U953 (N4637,N3933);
buff U954 (N4640,N3927);
buff U955 (N4643,N3948);
nor U956 (N4646,N490,N3948);
buff U957 (N4649,N3927);
buff U958 (N4652,N3933);
buff U959 (N4655,N3921);
buff U960 (N4658,N3942);
buff U961 (N4662,N3956);
buff U962 (N4665,N3948);
buff U963 (N4668,N3968);
buff U964 (N4671,N3962);
buff U965 (N4674,N3873);
buff U966 (N4677,N3867);
buff U967 (N4680,N3887);
buff U968 (N4683,N3881);
buff U969 (N4686,N3893);
buff U970 (N4689,N3849);
buff U971 (N4692,N3842);
buff U972 (N4695,N3861);
buff U973 (N4698,N3855);
nand U974 (N4701,N3813,N4223);
nand U975 (N4702,N3810,N4224);
not U976 (N4720,N4021);
nand U977 (N4721,N4021,N4263);
not U978 (N4724,N4147);
not U979 (N4725,N4144);
not U980 (N4726,N4159);
not U981 (N4727,N4156);
not U982 (N4728,N4153);
not U983 (N4729,N4097);
not U984 (N4730,N4094);
not U985 (N4731,N4091);
not U986 (N4732,N4088);
not U987 (N4733,N4109);
not U988 (N4734,N4106);
not U989 (N4735,N4103);
not U990 (N4736,N4100);
and U991 (N4737,N4273,N2877);
and U992 (N4738,N4274,N2877);
and U993 (N4739,N4276,N2877);
and U994 (N4740,N4277,N2877);
and U995 (N4741,N4150,N1758,N1755);
not U996 (N4855,N4212);
nand U997 (N4856,N4212,N2712);
nand U998 (N4908,N4215,N2718);
not U999 (N4909,N4215);
and U1000 (N4939,N4515,N4185);
and U1001 (N4942,N4516,N4186);
not U1002 (N4947,N4219);
and U1003 (N4953,N4188,N3775,N3779);
and U1004 (N4954,N3771,N4191,N3780);
and U1005 (N4955,N4191,N4188,N3038);
and U1006 (N4956,N4109,N3097,N3108);
and U1007 (N4957,N4106,N3097,N3108);
and U1008 (N4958,N4103,N3097,N3108);
and U1009 (N4959,N4100,N3097,N3108);
and U1010 (N4960,N4159,N3119,N3130);
and U1011 (N4961,N4156,N3119,N3130);
not U1012 (N4965,N4225);
not U1013 (N4966,N4228);
not U1014 (N4967,N4231);
not U1015 (N4968,N4234);
not U1016 (N4972,N4246);
not U1017 (N4973,N4249);
not U1018 (N4974,N4252);
nand U1019 (N4975,N4252,N4199);
not U1020 (N4976,N4206);
not U1021 (N4977,N4209);
and U1022 (N4978,N3793,N3789,N4206);
and U1023 (N4979,N4203,N4200,N4209);
and U1024 (N4980,N4097,N3147,N3158);
and U1025 (N4981,N4094,N3147,N3158);
and U1026 (N4982,N4091,N3147,N3158);
and U1027 (N4983,N4088,N3147,N3158);
and U1028 (N4984,N4153,N3169,N3180);
and U1029 (N4985,N4147,N3169,N3180);
and U1030 (N4986,N4144,N3169,N3180);
and U1031 (N4987,N4150,N3169,N3180);
nand U1032 (N5049,N4701,N4702);
not U1033 (N5052,N4237);
not U1034 (N5053,N4240);
not U1035 (N5054,N4243);
not U1036 (N5055,N4255);
not U1037 (N5056,N4258);
nand U1038 (N5057,N3819,N4720);
not U1039 (N5058,N4264);
nand U1040 (N5059,N4264,N4267);
and U1041 (N5060,N4724,N4725,N4269,N4027);
and U1042 (N5061,N4726,N4727,N3827,N4728);
and U1043 (N5062,N4729,N4730,N4731,N4732);
and U1044 (N5063,N4733,N4734,N4735,N4736);
and U1045 (N5065,N4357,N4375);
and U1046 (N5066,N4364,N4357,N4379);
and U1047 (N5067,N4418,N4436);
and U1048 (N5068,N4425,N4418,N4440);
not U1049 (N5069,N4548);
nand U1050 (N5070,N4548,N2628);
not U1051 (N5071,N4551);
nand U1052 (N5072,N4551,N2629);
not U1053 (N5073,N4554);
nand U1054 (N5074,N4554,N2630);
not U1055 (N5075,N4557);
nand U1056 (N5076,N4557,N2631);
not U1057 (N5077,N4560);
nand U1058 (N5078,N4560,N2632);
not U1059 (N5079,N4563);
nand U1060 (N5080,N4563,N2633);
not U1061 (N5081,N4566);
nand U1062 (N5082,N4566,N2634);
not U1063 (N5083,N4569);
nand U1064 (N5084,N4569,N2635);
not U1065 (N5085,N4572);
nand U1066 (N5086,N4572,N2636);
not U1067 (N5087,N4575);
nand U1068 (N5088,N4578,N2638);
not U1069 (N5089,N4578);
nand U1070 (N5090,N4581,N2639);
not U1071 (N5091,N4581);
nand U1072 (N5092,N4584,N2640);
not U1073 (N5093,N4584);
nand U1074 (N5094,N4587,N2641);
not U1075 (N5095,N4587);
nand U1076 (N5096,N4590,N2642);
not U1077 (N5097,N4590);
nand U1078 (N5098,N4593,N2643);
not U1079 (N5099,N4593);
nand U1080 (N5100,N4596,N2644);
not U1081 (N5101,N4596);
nand U1082 (N5102,N4599,N2645);
not U1083 (N5103,N4599);
nand U1084 (N5104,N4602,N2646);
not U1085 (N5105,N4602);
not U1086 (N5106,N4611);
nand U1087 (N5107,N4611,N2709);
not U1088 (N5108,N4614);
nand U1089 (N5109,N4614,N2710);
not U1090 (N5110,N4617);
nand U1091 (N5111,N4617,N2711);
nand U1092 (N5112,N1890,N4855);
not U1093 (N5113,N4621);
nand U1094 (N5114,N4621,N2713);
not U1095 (N5115,N4624);
nand U1096 (N5116,N4624,N2714);
and U1097 (N5117,N4364,N4379);
and U1098 (N5118,N4364,N4379);
and U1099 (N5119,N54,N4405);
not U1100 (N5120,N4627);
nand U1101 (N5121,N4630,N2716);
not U1102 (N5122,N4630);
nand U1103 (N5123,N4633,N2717);
not U1104 (N5124,N4633);
nand U1105 (N5125,N1908,N4909);
nand U1106 (N5126,N4637,N2719);
not U1107 (N5127,N4637);
nand U1108 (N5128,N4640,N2720);
not U1109 (N5129,N4640);
nand U1110 (N5130,N4643,N2721);
not U1111 (N5131,N4643);
and U1112 (N5132,N4425,N4440);
and U1113 (N5133,N4425,N4440);
not U1114 (N5135,N4649);
not U1115 (N5136,N4652);
nand U1116 (N5137,N4655,N4521);
not U1117 (N5138,N4655);
not U1118 (N5139,N4658);
nand U1119 (N5140,N4658,N4947);
not U1120 (N5141,N4674);
not U1121 (N5142,N4677);
not U1122 (N5143,N4680);
not U1123 (N5144,N4683);
nand U1124 (N5145,N4686,N4523);
not U1125 (N5146,N4686);
nor U1126 (N5147,N4953,N4196);
nor U1127 (N5148,N4954,N4955);
not U1128 (N5150,N4524);
nand U1129 (N5153,N4228,N4965);
nand U1130 (N5154,N4225,N4966);
nand U1131 (N5155,N4234,N4967);
nand U1132 (N5156,N4231,N4968);
not U1133 (N5157,N4532);
nand U1134 (N5160,N4249,N4972);
nand U1135 (N5161,N4246,N4973);
nand U1136 (N5162,N3816,N4974);
and U1137 (N5163,N4200,N3793,N4976);
and U1138 (N5164,N3789,N4203,N4977);
and U1139 (N5165,N4942,N3147,N3158);
not U1140 (N5166,N4512);
buff U1141 (N5169,N4290);
not U1142 (N5172,N4605);
buff U1143 (N5173,N4325);
not U1144 (N5176,N4608);
buff U1145 (N5177,N4349);
buff U1146 (N5180,N4405);
buff U1147 (N5183,N4357);
buff U1148 (N5186,N4357);
buff U1149 (N5189,N4364);
buff U1150 (N5192,N4364);
buff U1151 (N5195,N4385);
not U1152 (N5198,N4646);
buff U1153 (N5199,N4418);
buff U1154 (N5202,N4425);
buff U1155 (N5205,N4445);
buff U1156 (N5208,N4418);
buff U1157 (N5211,N4425);
buff U1158 (N5214,N4477);
buff U1159 (N5217,N4469);
buff U1160 (N5220,N4477);
not U1161 (N5223,N4662);
not U1162 (N5224,N4665);
not U1163 (N5225,N4668);
not U1164 (N5226,N4671);
not U1165 (N5227,N4689);
not U1166 (N5228,N4692);
not U1167 (N5229,N4695);
not U1168 (N5230,N4698);
nand U1169 (N5232,N4240,N5052);
nand U1170 (N5233,N4237,N5053);
nand U1171 (N5234,N4258,N5055);
nand U1172 (N5235,N4255,N5056);
nand U1173 (N5236,N4721,N5057);
nand U1174 (N5239,N3824,N5058);
and U1175 (N5240,N5060,N5061,N4270);
not U1176 (N5241,N4939);
nand U1177 (N5242,N1824,N5069);
nand U1178 (N5243,N1827,N5071);
nand U1179 (N5244,N1830,N5073);
nand U1180 (N5245,N1833,N5075);
nand U1181 (N5246,N1836,N5077);
nand U1182 (N5247,N1839,N5079);
nand U1183 (N5248,N1842,N5081);
nand U1184 (N5249,N1845,N5083);
nand U1185 (N5250,N1848,N5085);
nand U1186 (N5252,N1854,N5089);
nand U1187 (N5253,N1857,N5091);
nand U1188 (N5254,N1860,N5093);
nand U1189 (N5255,N1863,N5095);
nand U1190 (N5256,N1866,N5097);
nand U1191 (N5257,N1869,N5099);
nand U1192 (N5258,N1872,N5101);
nand U1193 (N5259,N1875,N5103);
nand U1194 (N5260,N1878,N5105);
nand U1195 (N5261,N1881,N5106);
nand U1196 (N5262,N1884,N5108);
nand U1197 (N5263,N1887,N5110);
nand U1198 (N5264,N5112,N4856);
nand U1199 (N5274,N1893,N5113);
nand U1200 (N5275,N1896,N5115);
nand U1201 (N5282,N1902,N5122);
nand U1202 (N5283,N1905,N5124);
nand U1203 (N5284,N4908,N5125);
nand U1204 (N5298,N1911,N5127);
nand U1205 (N5299,N1914,N5129);
nand U1206 (N5300,N1917,N5131);
nand U1207 (N5303,N4652,N5135);
nand U1208 (N5304,N4649,N5136);
nand U1209 (N5305,N4008,N5138);
nand U1210 (N5306,N4219,N5139);
nand U1211 (N5307,N4677,N5141);
nand U1212 (N5308,N4674,N5142);
nand U1213 (N5309,N4683,N5143);
nand U1214 (N5310,N4680,N5144);
nand U1215 (N5311,N4011,N5146);
not U1216 (N5312,N5049);
nand U1217 (N5315,N5153,N5154);
nand U1218 (N5319,N5155,N5156);
nand U1219 (N5324,N5160,N5161);
nand U1220 (N5328,N5162,N4975);
nor U1221 (N5331,N5163,N4978);
nor U1222 (N5332,N5164,N4979);
or U1223 (N5346,N4412,N5119);
nand U1224 (N5363,N4665,N5223);
nand U1225 (N5364,N4662,N5224);
nand U1226 (N5365,N4671,N5225);
nand U1227 (N5366,N4668,N5226);
nand U1228 (N5367,N4692,N5227);
nand U1229 (N5368,N4689,N5228);
nand U1230 (N5369,N4698,N5229);
nand U1231 (N5370,N4695,N5230);
nand U1232 (N5371,N5148,N5147);
buff U1233 (N5374,N4939);
nand U1234 (N5377,N5232,N5233);
nand U1235 (N5382,N5234,N5235);
nand U1236 (N5385,N5239,N5059);
and U1237 (N5388,N5062,N5063,N5241);
nand U1238 (N5389,N5242,N5070);
nand U1239 (N5396,N5243,N5072);
nand U1240 (N5407,N5244,N5074);
nand U1241 (N5418,N5245,N5076);
nand U1242 (N5424,N5246,N5078);
nand U1243 (N5431,N5247,N5080);
nand U1244 (N5441,N5248,N5082);
nand U1245 (N5452,N5249,N5084);
nand U1246 (N5462,N5250,N5086);
not U1247 (N5469,N5169);
nand U1248 (N5470,N5088,N5252);
nand U1249 (N5477,N5090,N5253);
nand U1250 (N5488,N5092,N5254);
nand U1251 (N5498,N5094,N5255);
nand U1252 (N5506,N5096,N5256);
nand U1253 (N5520,N5098,N5257);
nand U1254 (N5536,N5100,N5258);
nand U1255 (N5549,N5102,N5259);
nand U1256 (N5555,N5104,N5260);
nand U1257 (N5562,N5261,N5107);
nand U1258 (N5573,N5262,N5109);
nand U1259 (N5579,N5263,N5111);
nand U1260 (N5595,N5274,N5114);
nand U1261 (N5606,N5275,N5116);
nand U1262 (N5616,N5180,N2715);
not U1263 (N5617,N5180);
not U1264 (N5618,N5183);
not U1265 (N5619,N5186);
not U1266 (N5620,N5189);
not U1267 (N5621,N5192);
not U1268 (N5622,N5195);
nand U1269 (N5624,N5121,N5282);
nand U1270 (N5634,N5123,N5283);
nand U1271 (N5655,N5126,N5298);
nand U1272 (N5671,N5128,N5299);
nand U1273 (N5684,N5130,N5300);
not U1274 (N5690,N5202);
not U1275 (N5691,N5211);
nand U1276 (N5692,N5303,N5304);
nand U1277 (N5696,N5137,N5305);
nand U1278 (N5700,N5306,N5140);
nand U1279 (N5703,N5307,N5308);
nand U1280 (N5707,N5309,N5310);
nand U1281 (N5711,N5145,N5311);
and U1282 (N5726,N5166,N4512);
not U1283 (N5727,N5173);
not U1284 (N5728,N5177);
not U1285 (N5730,N5199);
not U1286 (N5731,N5205);
not U1287 (N5732,N5208);
not U1288 (N5733,N5214);
not U1289 (N5734,N5217);
not U1290 (N5735,N5220);
nand U1291 (N5736,N5365,N5366);
nand U1292 (N5739,N5363,N5364);
nand U1293 (N5742,N5369,N5370);
nand U1294 (N5745,N5367,N5368);
not U1295 (N5755,N5236);
nand U1296 (N5756,N5332,N5331);
and U1297 (N5954,N5264,N4396);
nand U1298 (N5955,N1899,N5617);
not U1299 (N5956,N5346);
and U1300 (N6005,N5284,N4456);
and U1301 (N6006,N5284,N4456);
not U1302 (N6023,N5371);
nand U1303 (N6024,N5371,N5312);
not U1304 (N6025,N5315);
not U1305 (N6028,N5324);
buff U1306 (N6031,N5319);
buff U1307 (N6034,N5319);
buff U1308 (N6037,N5328);
buff U1309 (N6040,N5328);
not U1310 (N6044,N5385);
or U1311 (N6045,N5166,N5726);
buff U1312 (N6048,N5264);
buff U1313 (N6051,N5284);
buff U1314 (N6054,N5284);
not U1315 (N6065,N5374);
nand U1316 (N6066,N5374,N5054);
not U1317 (N6067,N5377);
not U1318 (N6068,N5382);
nand U1319 (N6069,N5382,N5755);
and U1320 (N6071,N5470,N4316);
and U1321 (N6072,N5477,N5470,N4320);
and U1322 (N6073,N5488,N5470,N4325,N5477);
and U1323 (N6074,N5562,N4357,N4385,N4364);
and U1324 (N6075,N5389,N4280);
and U1325 (N6076,N5396,N5389,N4284);
and U1326 (N6077,N5407,N5389,N4290,N5396);
and U1327 (N6078,N5624,N4418,N4445,N4425);
not U1328 (N6079,N5418);
and U1329 (N6080,N5396,N5418,N5407,N5389);
and U1330 (N6083,N5396,N4284);
and U1331 (N6084,N5407,N4290,N5396);
and U1332 (N6085,N5418,N5407,N5396);
and U1333 (N6086,N5396,N4284);
and U1334 (N6087,N4290,N5407,N5396);
and U1335 (N6088,N5407,N4290);
and U1336 (N6089,N5418,N5407);
and U1337 (N6090,N5407,N4290);
and U1338 (N6091,N5431,N5462,N5441,N5424,N5452);
and U1339 (N6094,N5424,N4298);
and U1340 (N6095,N5431,N5424,N4301);
and U1341 (N6096,N5441,N5424,N4305,N5431);
and U1342 (N6097,N5452,N5441,N5424,N4310,N5431);
and U1343 (N6098,N5431,N4301);
and U1344 (N6099,N5441,N4305,N5431);
and U1345 (N6100,N5452,N5441,N4310,N5431);
and U1346 (N6101,N4,N5462,N5441,N5452,N5431);
and U1347 (N6102,N4305,N5441);
and U1348 (N6103,N5452,N5441,N4310);
and U1349 (N6104,N4,N5462,N5441,N5452);
and U1350 (N6105,N5452,N4310);
and U1351 (N6106,N4,N5462,N5452);
and U1352 (N6107,N4,N5462);
and U1353 (N6108,N5549,N5488,N5477,N5470);
and U1354 (N6111,N5477,N4320);
and U1355 (N6112,N5488,N4325,N5477);
and U1356 (N6113,N5549,N5488,N5477);
and U1357 (N6114,N5477,N4320);
and U1358 (N6115,N5488,N4325,N5477);
and U1359 (N6116,N5488,N4325);
and U1360 (N6117,N5555,N5536,N5520,N5506,N5498);
and U1361 (N6120,N5498,N4332);
and U1362 (N6121,N5506,N5498,N4336);
and U1363 (N6122,N5520,N5498,N4342,N5506);
and U1364 (N6123,N5536,N5520,N5498,N4349,N5506);
and U1365 (N6124,N5506,N4336);
and U1366 (N6125,N5520,N4342,N5506);
and U1367 (N6126,N5536,N5520,N4349,N5506);
and U1368 (N6127,N5555,N5520,N5506,N5536);
and U1369 (N6128,N5506,N4336);
and U1370 (N6129,N5520,N4342,N5506);
and U1371 (N6130,N5536,N5520,N4349,N5506);
and U1372 (N6131,N5520,N4342);
and U1373 (N6132,N5536,N5520,N4349);
and U1374 (N6133,N5555,N5520,N5536);
and U1375 (N6134,N5520,N4342);
and U1376 (N6135,N5536,N5520,N4349);
and U1377 (N6136,N5536,N4349);
and U1378 (N6137,N5549,N5488);
and U1379 (N6138,N5555,N5536);
not U1380 (N6139,N5573);
and U1381 (N6140,N4364,N5573,N5562,N4357);
and U1382 (N6143,N5562,N4385,N4364);
and U1383 (N6144,N5573,N5562,N4364);
and U1384 (N6145,N4385,N5562,N4364);
and U1385 (N6146,N5562,N4385);
and U1386 (N6147,N5573,N5562);
and U1387 (N6148,N5562,N4385);
and U1388 (N6149,N5264,N4405,N5595,N5579,N5606);
and U1389 (N6152,N5579,N4067);
and U1390 (N6153,N5264,N5579,N4396);
and U1391 (N6154,N5595,N5579,N4400,N5264);
and U1392 (N6155,N5606,N5595,N5579,N4412,N5264);
and U1393 (N6156,N5595,N4400,N5264);
and U1394 (N6157,N5606,N5595,N4412,N5264);
and U1395 (N6158,N54,N4405,N5595,N5606,N5264);
and U1396 (N6159,N4400,N5595);
and U1397 (N6160,N5606,N5595,N4412);
and U1398 (N6161,N54,N4405,N5595,N5606);
and U1399 (N6162,N5606,N4412);
and U1400 (N6163,N54,N4405,N5606);
nand U1401 (N6164,N5616,N5955);
and U1402 (N6168,N5684,N5624,N4425,N4418);
and U1403 (N6171,N5624,N4445,N4425);
and U1404 (N6172,N5684,N5624,N4425);
and U1405 (N6173,N5624,N4445,N4425);
and U1406 (N6174,N5624,N4445);
and U1407 (N6175,N4477,N5671,N5655,N5284,N5634);
and U1408 (N6178,N5634,N4080);
and U1409 (N6179,N5284,N5634,N4456);
and U1410 (N6180,N5655,N5634,N4462,N5284);
and U1411 (N6181,N5671,N5655,N5634,N4469,N5284);
and U1412 (N6182,N5655,N4462,N5284);
and U1413 (N6183,N5671,N5655,N4469,N5284);
and U1414 (N6184,N4477,N5655,N5284,N5671);
and U1415 (N6185,N5655,N4462,N5284);
and U1416 (N6186,N5671,N5655,N4469,N5284);
and U1417 (N6187,N5655,N4462);
and U1418 (N6188,N5671,N5655,N4469);
and U1419 (N6189,N4477,N5655,N5671);
and U1420 (N6190,N5655,N4462);
and U1421 (N6191,N5671,N5655,N4469);
and U1422 (N6192,N5671,N4469);
and U1423 (N6193,N5684,N5624);
and U1424 (N6194,N4477,N5671);
not U1425 (N6197,N5692);
not U1426 (N6200,N5696);
not U1427 (N6203,N5703);
not U1428 (N6206,N5707);
buff U1429 (N6209,N5700);
buff U1430 (N6212,N5700);
buff U1431 (N6215,N5711);
buff U1432 (N6218,N5711);
nand U1433 (N6221,N5049,N6023);
not U1434 (N6234,N5756);
nand U1435 (N6235,N5756,N6044);
buff U1436 (N6238,N5462);
buff U1437 (N6241,N5389);
buff U1438 (N6244,N5389);
buff U1439 (N6247,N5396);
buff U1440 (N6250,N5396);
buff U1441 (N6253,N5407);
buff U1442 (N6256,N5407);
buff U1443 (N6259,N5424);
buff U1444 (N6262,N5431);
buff U1445 (N6265,N5441);
buff U1446 (N6268,N5452);
buff U1447 (N6271,N5549);
buff U1448 (N6274,N5488);
buff U1449 (N6277,N5470);
buff U1450 (N6280,N5477);
buff U1451 (N6283,N5549);
buff U1452 (N6286,N5488);
buff U1453 (N6289,N5470);
buff U1454 (N6292,N5477);
buff U1455 (N6295,N5555);
buff U1456 (N6298,N5536);
buff U1457 (N6301,N5498);
buff U1458 (N6304,N5520);
buff U1459 (N6307,N5506);
buff U1460 (N6310,N5506);
buff U1461 (N6313,N5555);
buff U1462 (N6316,N5536);
buff U1463 (N6319,N5498);
buff U1464 (N6322,N5520);
buff U1465 (N6325,N5562);
buff U1466 (N6328,N5562);
buff U1467 (N6331,N5579);
buff U1468 (N6335,N5595);
buff U1469 (N6338,N5606);
buff U1470 (N6341,N5684);
buff U1471 (N6344,N5624);
buff U1472 (N6347,N5684);
buff U1473 (N6350,N5624);
buff U1474 (N6353,N5671);
buff U1475 (N6356,N5634);
buff U1476 (N6359,N5655);
buff U1477 (N6364,N5671);
buff U1478 (N6367,N5634);
buff U1479 (N6370,N5655);
not U1480 (N6373,N5736);
not U1481 (N6374,N5739);
not U1482 (N6375,N5742);
not U1483 (N6376,N5745);
nand U1484 (N6377,N4243,N6065);
nand U1485 (N6378,N5236,N6068);
or U1486 (N6382,N4268,N6071,N6072,N6073);
or U1487 (N6386,N3968,N5065,N5066,N6074);
or U1488 (N6388,N4271,N6075,N6076,N6077);
or U1489 (N6392,N3968,N5067,N5068,N6078);
or U1490 (N6397,N4297,N6094,N6095,N6096,N6097);
or U1491 (N6411,N4320,N6116);
or U1492 (N6415,N4331,N6120,N6121,N6122,N6123);
or U1493 (N6419,N4342,N6136);
or U1494 (N6427,N4392,N6152,N6153,N6154,N6155);
not U1495 (N6434,N6048);
or U1496 (N6437,N4440,N6174);
or U1497 (N6441,N4451,N6178,N6179,N6180,N6181);
or U1498 (N6445,N4462,N6192);
not U1499 (N6448,N6051);
not U1500 (N6449,N6054);
nand U1501 (N6466,N6221,N6024);
not U1502 (N6469,N6031);
not U1503 (N6470,N6034);
not U1504 (N6471,N6037);
not U1505 (N6472,N6040);
and U1506 (N6473,N5315,N4524,N6031);
and U1507 (N6474,N6025,N5150,N6034);
and U1508 (N6475,N5324,N4532,N6037);
and U1509 (N6476,N6028,N5157,N6040);
nand U1510 (N6477,N5385,N6234);
nand U1511 (N6478,N6045,N132);
or U1512 (N6482,N4280,N6083,N6084,N6085);
nor U1513 (N6486,N4280,N6086,N6087);
or U1514 (N6490,N4284,N6088,N6089);
nor U1515 (N6494,N4284,N6090);
or U1516 (N6500,N4298,N6098,N6099,N6100,N6101);
or U1517 (N6504,N4301,N6102,N6103,N6104);
or U1518 (N6508,N4305,N6105,N6106);
or U1519 (N6512,N4310,N6107);
or U1520 (N6516,N4316,N6111,N6112,N6113);
nor U1521 (N6526,N4316,N6114,N6115);
or U1522 (N6536,N4336,N6131,N6132,N6133);
or U1523 (N6539,N4332,N6124,N6125,N6126,N6127);
nor U1524 (N6553,N4336,N6134,N6135);
nor U1525 (N6556,N4332,N6128,N6129,N6130);
or U1526 (N6566,N4375,N5117,N6143,N6144);
nor U1527 (N6569,N4375,N5118,N6145);
or U1528 (N6572,N4379,N6146,N6147);
nor U1529 (N6575,N4379,N6148);
or U1530 (N6580,N4067,N5954,N6156,N6157,N6158);
or U1531 (N6584,N4396,N6159,N6160,N6161);
or U1532 (N6587,N4400,N6162,N6163);
or U1533 (N6592,N4436,N5132,N6171,N6172);
nor U1534 (N6599,N4436,N5133,N6173);
or U1535 (N6606,N4456,N6187,N6188,N6189);
or U1536 (N6609,N4080,N6005,N6182,N6183,N6184);
nor U1537 (N6619,N4456,N6190,N6191);
nor U1538 (N6622,N4080,N6006,N6185,N6186);
nand U1539 (N6630,N5739,N6373);
nand U1540 (N6631,N5736,N6374);
nand U1541 (N6632,N5745,N6375);
nand U1542 (N6633,N5742,N6376);
nand U1543 (N6634,N6377,N6066);
nand U1544 (N6637,N6069,N6378);
not U1545 (N6640,N6164);
and U1546 (N6641,N6108,N6117);
and U1547 (N6643,N6140,N6149);
and U1548 (N6646,N6168,N6175);
and U1549 (N6648,N6080,N6091);
nand U1550 (N6650,N6238,N2637);
not U1551 (N6651,N6238);
not U1552 (N6653,N6241);
not U1553 (N6655,N6244);
not U1554 (N6657,N6247);
not U1555 (N6659,N6250);
nand U1556 (N6660,N6253,N5087);
not U1557 (N6661,N6253);
nand U1558 (N6662,N6256,N5469);
not U1559 (N6663,N6256);
and U1560 (N6664,N6091,N4);
not U1561 (N6666,N6259);
not U1562 (N6668,N6262);
not U1563 (N6670,N6265);
not U1564 (N6672,N6268);
not U1565 (N6675,N6117);
not U1566 (N6680,N6280);
not U1567 (N6681,N6292);
not U1568 (N6682,N6307);
not U1569 (N6683,N6310);
nand U1570 (N6689,N6325,N5120);
not U1571 (N6690,N6325);
nand U1572 (N6691,N6328,N5622);
not U1573 (N6692,N6328);
and U1574 (N6693,N6149,N54);
not U1575 (N6695,N6331);
not U1576 (N6698,N6335);
nand U1577 (N6699,N6338,N5956);
not U1578 (N6700,N6338);
not U1579 (N6703,N6175);
not U1580 (N6708,N6209);
not U1581 (N6709,N6212);
not U1582 (N6710,N6215);
not U1583 (N6711,N6218);
and U1584 (N6712,N5696,N5692,N6209);
and U1585 (N6713,N6200,N6197,N6212);
and U1586 (N6714,N5707,N5703,N6215);
and U1587 (N6715,N6206,N6203,N6218);
buff U1588 (N6716,N6466);
and U1589 (N6718,N6164,N1777,N3130);
and U1590 (N6719,N5150,N5315,N6469);
and U1591 (N6720,N4524,N6025,N6470);
and U1592 (N6721,N5157,N5324,N6471);
and U1593 (N6722,N4532,N6028,N6472);
nand U1594 (N6724,N6477,N6235);
not U1595 (N6739,N6271);
not U1596 (N6740,N6274);
not U1597 (N6741,N6277);
not U1598 (N6744,N6283);
not U1599 (N6745,N6286);
not U1600 (N6746,N6289);
not U1601 (N6751,N6295);
not U1602 (N6752,N6298);
not U1603 (N6753,N6301);
not U1604 (N6754,N6304);
not U1605 (N6755,N6322);
not U1606 (N6760,N6313);
not U1607 (N6761,N6316);
not U1608 (N6762,N6319);
not U1609 (N6772,N6341);
not U1610 (N6773,N6344);
not U1611 (N6776,N6347);
not U1612 (N6777,N6350);
not U1613 (N6782,N6353);
not U1614 (N6783,N6356);
not U1615 (N6784,N6359);
not U1616 (N6785,N6370);
not U1617 (N6790,N6364);
not U1618 (N6791,N6367);
nand U1619 (N6792,N6630,N6631);
nand U1620 (N6795,N6632,N6633);
and U1621 (N6801,N6108,N6415);
and U1622 (N6802,N6427,N6140);
and U1623 (N6803,N6397,N6080);
and U1624 (N6804,N6168,N6441);
not U1625 (N6805,N6466);
nand U1626 (N6806,N1851,N6651);
not U1627 (N6807,N6482);
nand U1628 (N6808,N6482,N6653);
not U1629 (N6809,N6486);
nand U1630 (N6810,N6486,N6655);
not U1631 (N6811,N6490);
nand U1632 (N6812,N6490,N6657);
not U1633 (N6813,N6494);
nand U1634 (N6814,N6494,N6659);
nand U1635 (N6815,N4575,N6661);
nand U1636 (N6816,N5169,N6663);
or U1637 (N6817,N6397,N6664);
not U1638 (N6823,N6500);
nand U1639 (N6824,N6500,N6666);
not U1640 (N6825,N6504);
nand U1641 (N6826,N6504,N6668);
not U1642 (N6827,N6508);
nand U1643 (N6828,N6508,N6670);
not U1644 (N6829,N6512);
nand U1645 (N6830,N6512,N6672);
not U1646 (N6831,N6415);
not U1647 (N6834,N6566);
nand U1648 (N6835,N6566,N5618);
not U1649 (N6836,N6569);
nand U1650 (N6837,N6569,N5619);
not U1651 (N6838,N6572);
nand U1652 (N6839,N6572,N5620);
not U1653 (N6840,N6575);
nand U1654 (N6841,N6575,N5621);
nand U1655 (N6842,N4627,N6690);
nand U1656 (N6843,N5195,N6692);
or U1657 (N6844,N6427,N6693);
not U1658 (N6850,N6580);
nand U1659 (N6851,N6580,N6695);
not U1660 (N6852,N6584);
nand U1661 (N6853,N6584,N6434);
not U1662 (N6854,N6587);
nand U1663 (N6855,N6587,N6698);
nand U1664 (N6856,N5346,N6700);
not U1665 (N6857,N6441);
and U1666 (N6860,N6197,N5696,N6708);
and U1667 (N6861,N5692,N6200,N6709);
and U1668 (N6862,N6203,N5707,N6710);
and U1669 (N6863,N5703,N6206,N6711);
or U1670 (N6866,N4197,N6718,N3785);
nor U1671 (N6872,N6719,N6473);
nor U1672 (N6873,N6720,N6474);
nor U1673 (N6874,N6721,N6475);
nor U1674 (N6875,N6722,N6476);
not U1675 (N6876,N6637);
buff U1676 (N6877,N6724);
and U1677 (N6879,N6045,N6478);
and U1678 (N6880,N6478,N132);
or U1679 (N6881,N6411,N6137);
not U1680 (N6884,N6516);
not U1681 (N6885,N6411);
not U1682 (N6888,N6526);
not U1683 (N6889,N6536);
nand U1684 (N6890,N6536,N5176);
or U1685 (N6891,N6419,N6138);
not U1686 (N6894,N6539);
not U1687 (N6895,N6553);
nand U1688 (N6896,N6553,N5728);
not U1689 (N6897,N6419);
not U1690 (N6900,N6556);
or U1691 (N6901,N6437,N6193);
not U1692 (N6904,N6592);
not U1693 (N6905,N6437);
not U1694 (N6908,N6599);
or U1695 (N6909,N6445,N6194);
not U1696 (N6912,N6606);
not U1697 (N6913,N6609);
not U1698 (N6914,N6619);
nand U1699 (N6915,N6619,N5734);
not U1700 (N6916,N6445);
not U1701 (N6919,N6622);
not U1702 (N6922,N6634);
nand U1703 (N6923,N6634,N6067);
or U1704 (N6924,N6382,N6801);
or U1705 (N6925,N6386,N6802);
or U1706 (N6926,N6388,N6803);
or U1707 (N6927,N6392,N6804);
not U1708 (N6930,N6724);
nand U1709 (N6932,N6650,N6806);
nand U1710 (N6935,N6241,N6807);
nand U1711 (N6936,N6244,N6809);
nand U1712 (N6937,N6247,N6811);
nand U1713 (N6938,N6250,N6813);
nand U1714 (N6939,N6660,N6815);
nand U1715 (N6940,N6662,N6816);
nand U1716 (N6946,N6259,N6823);
nand U1717 (N6947,N6262,N6825);
nand U1718 (N6948,N6265,N6827);
nand U1719 (N6949,N6268,N6829);
nand U1720 (N6953,N5183,N6834);
nand U1721 (N6954,N5186,N6836);
nand U1722 (N6955,N5189,N6838);
nand U1723 (N6956,N5192,N6840);
nand U1724 (N6957,N6689,N6842);
nand U1725 (N6958,N6691,N6843);
nand U1726 (N6964,N6331,N6850);
nand U1727 (N6965,N6048,N6852);
nand U1728 (N6966,N6335,N6854);
nand U1729 (N6967,N6699,N6856);
nor U1730 (N6973,N6860,N6712);
nor U1731 (N6974,N6861,N6713);
nor U1732 (N6975,N6862,N6714);
nor U1733 (N6976,N6863,N6715);
not U1734 (N6977,N6792);
not U1735 (N6978,N6795);
or U1736 (N6979,N6879,N6880);
nand U1737 (N6987,N4608,N6889);
nand U1738 (N6990,N5177,N6895);
nand U1739 (N6999,N5217,N6914);
nand U1740 (N7002,N5377,N6922);
nand U1741 (N7003,N6873,N6872);
nand U1742 (N7006,N6875,N6874);
and U1743 (N7011,N6866,N2681,N2692);
and U1744 (N7012,N6866,N2756,N2767);
and U1745 (N7013,N6866,N2779,N2790);
not U1746 (N7015,N6866);
and U1747 (N7016,N6866,N2801,N2812);
nand U1748 (N7018,N6935,N6808);
nand U1749 (N7019,N6936,N6810);
nand U1750 (N7020,N6937,N6812);
nand U1751 (N7021,N6938,N6814);
not U1752 (N7022,N6939);
not U1753 (N7023,N6817);
nand U1754 (N7028,N6946,N6824);
nand U1755 (N7031,N6947,N6826);
nand U1756 (N7034,N6948,N6828);
nand U1757 (N7037,N6949,N6830);
and U1758 (N7040,N6817,N6079);
and U1759 (N7041,N6831,N6675);
nand U1760 (N7044,N6953,N6835);
nand U1761 (N7045,N6954,N6837);
nand U1762 (N7046,N6955,N6839);
nand U1763 (N7047,N6956,N6841);
not U1764 (N7048,N6957);
not U1765 (N7049,N6844);
nand U1766 (N7054,N6964,N6851);
nand U1767 (N7057,N6965,N6853);
nand U1768 (N7060,N6966,N6855);
and U1769 (N7064,N6844,N6139);
and U1770 (N7065,N6857,N6703);
not U1771 (N7072,N6881);
nand U1772 (N7073,N6881,N5172);
not U1773 (N7074,N6885);
nand U1774 (N7075,N6885,N5727);
nand U1775 (N7076,N6890,N6987);
not U1776 (N7079,N6891);
nand U1777 (N7080,N6896,N6990);
not U1778 (N7083,N6897);
not U1779 (N7084,N6901);
nand U1780 (N7085,N6901,N5198);
not U1781 (N7086,N6905);
nand U1782 (N7087,N6905,N5731);
not U1783 (N7088,N6909);
nand U1784 (N7089,N6909,N6912);
nand U1785 (N7090,N6915,N6999);
not U1786 (N7093,N6916);
nand U1787 (N7094,N6974,N6973);
nand U1788 (N7097,N6976,N6975);
nand U1789 (N7101,N7002,N6923);
not U1790 (N7105,N6932);
not U1791 (N7110,N6967);
and U1792 (N7114,N6979,N603,N1755);
not U1793 (N7115,N7019);
not U1794 (N7116,N7021);
and U1795 (N7125,N6817,N7018);
and U1796 (N7126,N6817,N7020);
and U1797 (N7127,N6817,N7022);
not U1798 (N7130,N7045);
not U1799 (N7131,N7047);
and U1800 (N7139,N6844,N7044);
and U1801 (N7140,N6844,N7046);
and U1802 (N7141,N6844,N7048);
and U1803 (N7146,N6932,N1761,N3108);
and U1804 (N7147,N6967,N1777,N3130);
not U1805 (N7149,N7003);
not U1806 (N7150,N7006);
nand U1807 (N7151,N7006,N6876);
nand U1808 (N7152,N4605,N7072);
nand U1809 (N7153,N5173,N7074);
nand U1810 (N7158,N4646,N7084);
nand U1811 (N7159,N5205,N7086);
nand U1812 (N7160,N6606,N7088);
not U1813 (N7166,N7037);
not U1814 (N7167,N7034);
not U1815 (N7168,N7031);
not U1816 (N7169,N7028);
not U1817 (N7170,N7060);
not U1818 (N7171,N7057);
not U1819 (N7172,N7054);
and U1820 (N7173,N7115,N7023);
and U1821 (N7174,N7116,N7023);
and U1822 (N7175,N6940,N7023);
and U1823 (N7176,N5418,N7023);
not U1824 (N7177,N7041);
and U1825 (N7178,N7130,N7049);
and U1826 (N7179,N7131,N7049);
and U1827 (N7180,N6958,N7049);
and U1828 (N7181,N5573,N7049);
not U1829 (N7182,N7065);
not U1830 (N7183,N7094);
nand U1831 (N7184,N7094,N6977);
not U1832 (N7185,N7097);
nand U1833 (N7186,N7097,N6978);
and U1834 (N7187,N7037,N1761,N3108);
and U1835 (N7188,N7034,N1761,N3108);
and U1836 (N7189,N7031,N1761,N3108);
or U1837 (N7190,N4956,N7146,N3781);
and U1838 (N7196,N7060,N1777,N3130);
and U1839 (N7197,N7057,N1777,N3130);
or U1840 (N7198,N4960,N7147,N3786);
nand U1841 (N7204,N7101,N7149);
not U1842 (N7205,N7101);
nand U1843 (N7206,N6637,N7150);
and U1844 (N7207,N7028,N1793,N3158);
and U1845 (N7208,N7054,N1807,N3180);
nand U1846 (N7209,N7073,N7152);
nand U1847 (N7212,N7075,N7153);
not U1848 (N7215,N7076);
nand U1849 (N7216,N7076,N7079);
not U1850 (N7217,N7080);
nand U1851 (N7218,N7080,N7083);
nand U1852 (N7219,N7085,N7158);
nand U1853 (N7222,N7087,N7159);
nand U1854 (N7225,N7089,N7160);
not U1855 (N7228,N7090);
nand U1856 (N7229,N7090,N7093);
or U1857 (N7236,N7173,N7125);
or U1858 (N7239,N7174,N7126);
or U1859 (N7242,N7175,N7127);
or U1860 (N7245,N7176,N7040);
or U1861 (N7250,N7178,N7139);
or U1862 (N7257,N7179,N7140);
or U1863 (N7260,N7180,N7141);
or U1864 (N7263,N7181,N7064);
nand U1865 (N7268,N6792,N7183);
nand U1866 (N7269,N6795,N7185);
or U1867 (N7270,N4957,N7187,N3782);
or U1868 (N7276,N4958,N7188,N3783);
or U1869 (N7282,N4959,N7189,N3784);
or U1870 (N7288,N4961,N7196,N3787);
or U1871 (N7294,N3998,N7197,N3788);
nand U1872 (N7300,N7003,N7205);
nand U1873 (N7301,N7206,N7151);
or U1874 (N7304,N4980,N7207,N3800);
or U1875 (N7310,N4984,N7208,N3805);
nand U1876 (N7320,N6891,N7215);
nand U1877 (N7321,N6897,N7217);
nand U1878 (N7328,N6916,N7228);
and U1879 (N7338,N7190,N1185,N2692);
and U1880 (N7339,N7198,N2681,N2692);
and U1881 (N7340,N7190,N1247,N2767);
and U1882 (N7341,N7198,N2756,N2767);
and U1883 (N7342,N7190,N1327,N2790);
and U1884 (N7349,N7198,N2779,N2790);
and U1885 (N7357,N7198,N2801,N2812);
not U1886 (N7363,N7198);
and U1887 (N7364,N7190,N1351,N2812);
not U1888 (N7365,N7190);
nand U1889 (N7394,N7268,N7184);
nand U1890 (N7397,N7269,N7186);
nand U1891 (N7402,N7204,N7300);
not U1892 (N7405,N7209);
nand U1893 (N7406,N7209,N6884);
not U1894 (N7407,N7212);
nand U1895 (N7408,N7212,N6888);
nand U1896 (N7409,N7320,N7216);
nand U1897 (N7412,N7321,N7218);
not U1898 (N7415,N7219);
nand U1899 (N7416,N7219,N6904);
not U1900 (N7417,N7222);
nand U1901 (N7418,N7222,N6908);
not U1902 (N7419,N7225);
nand U1903 (N7420,N7225,N6913);
nand U1904 (N7421,N7328,N7229);
not U1905 (N7424,N7245);
not U1906 (N7425,N7242);
not U1907 (N7426,N7239);
not U1908 (N7427,N7236);
not U1909 (N7428,N7263);
not U1910 (N7429,N7260);
not U1911 (N7430,N7257);
not U1912 (N7431,N7250);
not U1913 (N7432,N7250);
and U1914 (N7433,N7310,N2653,N2664);
and U1915 (N7434,N7304,N1161,N2664);
or U1916 (N7435,N7011,N7338,N3621,N2591);
and U1917 (N7436,N7270,N1185,N2692);
and U1918 (N7437,N7288,N2681,N2692);
and U1919 (N7438,N7276,N1185,N2692);
and U1920 (N7439,N7294,N2681,N2692);
and U1921 (N7440,N7282,N1185,N2692);
and U1922 (N7441,N7310,N2728,N2739);
and U1923 (N7442,N7304,N1223,N2739);
or U1924 (N7443,N7012,N7340,N3632,N2600);
and U1925 (N7444,N7270,N1247,N2767);
and U1926 (N7445,N7288,N2756,N2767);
and U1927 (N7446,N7276,N1247,N2767);
and U1928 (N7447,N7294,N2756,N2767);
and U1929 (N7448,N7282,N1247,N2767);
or U1930 (N7449,N7013,N7342,N3641,N2605);
and U1931 (N7450,N7310,N3041,N3052);
and U1932 (N7451,N7304,N1697,N3052);
and U1933 (N7452,N7294,N2779,N2790);
and U1934 (N7453,N7282,N1327,N2790);
and U1935 (N7454,N7288,N2779,N2790);
and U1936 (N7455,N7276,N1327,N2790);
and U1937 (N7456,N7270,N1327,N2790);
and U1938 (N7457,N7310,N3075,N3086);
and U1939 (N7458,N7304,N1731,N3086);
and U1940 (N7459,N7294,N2801,N2812);
and U1941 (N7460,N7282,N1351,N2812);
and U1942 (N7461,N7288,N2801,N2812);
and U1943 (N7462,N7276,N1351,N2812);
and U1944 (N7463,N7270,N1351,N2812);
and U1945 (N7464,N7250,N603,N599);
not U1946 (N7465,N7310);
not U1947 (N7466,N7294);
not U1948 (N7467,N7288);
not U1949 (N7468,N7301);
or U1950 (N7469,N7016,N7364,N3660,N2626);
not U1951 (N7470,N7304);
not U1952 (N7471,N7282);
not U1953 (N7472,N7276);
not U1954 (N7473,N7270);
buff U1955 (N7474,N7394);
buff U1956 (N7476,N7397);
and U1957 (N7479,N7301,N3068);
and U1958 (N7481,N7245,N1793,N3158);
and U1959 (N7482,N7242,N1793,N3158);
and U1960 (N7483,N7239,N1793,N3158);
and U1961 (N7484,N7236,N1793,N3158);
and U1962 (N7485,N7263,N1807,N3180);
and U1963 (N7486,N7260,N1807,N3180);
and U1964 (N7487,N7257,N1807,N3180);
and U1965 (N7488,N7250,N1807,N3180);
nand U1966 (N7489,N6979,N7250);
nand U1967 (N7492,N6516,N7405);
nand U1968 (N7493,N6526,N7407);
nand U1969 (N7498,N6592,N7415);
nand U1970 (N7499,N6599,N7417);
nand U1971 (N7500,N6609,N7419);
and U1972 (N7503,N7105,N7166,N7167,N7168,N7169,N7424,N7425,N7426,N7427);
and U1973 (N7504,N6640,N7110,N7170,N7171,N7172,N7428,N7429,N7430,N7431);
or U1974 (N7505,N7433,N7434,N3616,N2585);
and U1975 (N7506,N7435,N2675);
or U1976 (N7507,N7339,N7436,N3622,N2592);
or U1977 (N7508,N7437,N7438,N3623,N2593);
or U1978 (N7509,N7439,N7440,N3624,N2594);
or U1979 (N7510,N7441,N7442,N3627,N2595);
and U1980 (N7511,N7443,N2750);
or U1981 (N7512,N7341,N7444,N3633,N2601);
or U1982 (N7513,N7445,N7446,N3634,N2602);
or U1983 (N7514,N7447,N7448,N3635,N2603);
or U1984 (N7515,N7450,N7451,N3646,N2610);
or U1985 (N7516,N7452,N7453,N3647,N2611);
or U1986 (N7517,N7454,N7455,N3648,N2612);
or U1987 (N7518,N7349,N7456,N3649,N2613);
or U1988 (N7519,N7457,N7458,N3654,N2618);
or U1989 (N7520,N7459,N7460,N3655,N2619);
or U1990 (N7521,N7461,N7462,N3656,N2620);
or U1991 (N7522,N7357,N7463,N3657,N2621);
or U1992 (N7525,N4741,N7114,N2624,N7464);
and U1993 (N7526,N7468,N3119,N3130);
not U1994 (N7527,N7394);
not U1995 (N7528,N7397);
not U1996 (N7529,N7402);
and U1997 (N7530,N7402,N3068);
or U1998 (N7531,N4981,N7481,N3801);
or U1999 (N7537,N4982,N7482,N3802);
or U2000 (N7543,N4983,N7483,N3803);
or U2001 (N7549,N5165,N7484,N3804);
or U2002 (N7555,N4985,N7485,N3806);
or U2003 (N7561,N4986,N7486,N3807);
or U2004 (N7567,N4547,N7487,N3808);
or U2005 (N7573,N4987,N7488,N3809);
nand U2006 (N7579,N7492,N7406);
nand U2007 (N7582,N7493,N7408);
not U2008 (N7585,N7409);
nand U2009 (N7586,N7409,N6894);
not U2010 (N7587,N7412);
nand U2011 (N7588,N7412,N6900);
nand U2012 (N7589,N7498,N7416);
nand U2013 (N7592,N7499,N7418);
nand U2014 (N7595,N7500,N7420);
not U2015 (N7598,N7421);
nand U2016 (N7599,N7421,N6919);
and U2017 (N7600,N7505,N2647);
and U2018 (N7601,N7507,N2675);
and U2019 (N7602,N7508,N2675);
and U2020 (N7603,N7509,N2675);
and U2021 (N7604,N7510,N2722);
and U2022 (N7605,N7512,N2750);
and U2023 (N7606,N7513,N2750);
and U2024 (N7607,N7514,N2750);
and U2025 (N7624,N6979,N7489);
and U2026 (N7625,N7489,N7250);
and U2027 (N7626,N1149,N7525);
and U2028 (N7631,N562,N7527,N7528,N6805,N6930);
and U2029 (N7636,N7529,N3097,N3108);
nand U2030 (N7657,N6539,N7585);
nand U2031 (N7658,N6556,N7587);
nand U2032 (N7665,N6622,N7598);
and U2033 (N7666,N7555,N2653,N2664);
and U2034 (N7667,N7531,N1161,N2664);
and U2035 (N7668,N7561,N2653,N2664);
and U2036 (N7669,N7537,N1161,N2664);
and U2037 (N7670,N7567,N2653,N2664);
and U2038 (N7671,N7543,N1161,N2664);
and U2039 (N7672,N7573,N2653,N2664);
and U2040 (N7673,N7549,N1161,N2664);
and U2041 (N7674,N7555,N2728,N2739);
and U2042 (N7675,N7531,N1223,N2739);
and U2043 (N7676,N7561,N2728,N2739);
and U2044 (N7677,N7537,N1223,N2739);
and U2045 (N7678,N7567,N2728,N2739);
and U2046 (N7679,N7543,N1223,N2739);
and U2047 (N7680,N7573,N2728,N2739);
and U2048 (N7681,N7549,N1223,N2739);
and U2049 (N7682,N7573,N3075,N3086);
and U2050 (N7683,N7549,N1731,N3086);
and U2051 (N7684,N7573,N3041,N3052);
and U2052 (N7685,N7549,N1697,N3052);
and U2053 (N7686,N7567,N3041,N3052);
and U2054 (N7687,N7543,N1697,N3052);
and U2055 (N7688,N7561,N3041,N3052);
and U2056 (N7689,N7537,N1697,N3052);
and U2057 (N7690,N7555,N3041,N3052);
and U2058 (N7691,N7531,N1697,N3052);
and U2059 (N7692,N7567,N3075,N3086);
and U2060 (N7693,N7543,N1731,N3086);
and U2061 (N7694,N7561,N3075,N3086);
and U2062 (N7695,N7537,N1731,N3086);
and U2063 (N7696,N7555,N3075,N3086);
and U2064 (N7697,N7531,N1731,N3086);
or U2065 (N7698,N7624,N7625);
not U2066 (N7699,N7573);
not U2067 (N7700,N7567);
not U2068 (N7701,N7561);
not U2069 (N7702,N7555);
and U2070 (N7703,N1156,N7631,N245);
not U2071 (N7704,N7549);
not U2072 (N7705,N7543);
not U2073 (N7706,N7537);
not U2074 (N7707,N7531);
not U2075 (N7708,N7579);
nand U2076 (N7709,N7579,N6739);
not U2077 (N7710,N7582);
nand U2078 (N7711,N7582,N6744);
nand U2079 (N7712,N7657,N7586);
nand U2080 (N7715,N7658,N7588);
not U2081 (N7718,N7589);
nand U2082 (N7719,N7589,N6772);
not U2083 (N7720,N7592);
nand U2084 (N7721,N7592,N6776);
not U2085 (N7722,N7595);
nand U2086 (N7723,N7595,N5733);
nand U2087 (N7724,N7665,N7599);
or U2088 (N7727,N7666,N7667,N3617,N2586);
or U2089 (N7728,N7668,N7669,N3618,N2587);
or U2090 (N7729,N7670,N7671,N3619,N2588);
or U2091 (N7730,N7672,N7673,N3620,N2589);
or U2092 (N7731,N7674,N7675,N3628,N2596);
or U2093 (N7732,N7676,N7677,N3629,N2597);
or U2094 (N7733,N7678,N7679,N3630,N2598);
or U2095 (N7734,N7680,N7681,N3631,N2599);
or U2096 (N7735,N7682,N7683,N3638,N2604);
or U2097 (N7736,N7684,N7685,N3642,N2606);
or U2098 (N7737,N7686,N7687,N3643,N2607);
or U2099 (N7738,N7688,N7689,N3644,N2608);
or U2100 (N7739,N7690,N7691,N3645,N2609);
or U2101 (N7740,N7692,N7693,N3651,N2615);
or U2102 (N7741,N7694,N7695,N3652,N2616);
or U2103 (N7742,N7696,N7697,N3653,N2617);
nand U2104 (N7743,N6271,N7708);
nand U2105 (N7744,N6283,N7710);
nand U2106 (N7749,N6341,N7718);
nand U2107 (N7750,N6347,N7720);
nand U2108 (N7751,N5214,N7722);
and U2109 (N7754,N7727,N2647);
and U2110 (N7755,N7728,N2647);
and U2111 (N7756,N7729,N2647);
and U2112 (N7757,N7730,N2647);
and U2113 (N7758,N7731,N2722);
and U2114 (N7759,N7732,N2722);
and U2115 (N7760,N7733,N2722);
and U2116 (N7761,N7734,N2722);
nand U2117 (N7762,N7743,N7709);
nand U2118 (N7765,N7744,N7711);
not U2119 (N7768,N7712);
nand U2120 (N7769,N7712,N6751);
not U2121 (N7770,N7715);
nand U2122 (N7771,N7715,N6760);
nand U2123 (N7772,N7749,N7719);
nand U2124 (N7775,N7750,N7721);
nand U2125 (N7778,N7751,N7723);
not U2126 (N7781,N7724);
nand U2127 (N7782,N7724,N5735);
nand U2128 (N7787,N6295,N7768);
nand U2129 (N7788,N6313,N7770);
nand U2130 (N7795,N5220,N7781);
not U2131 (N7796,N7762);
nand U2132 (N7797,N7762,N6740);
not U2133 (N7798,N7765);
nand U2134 (N7799,N7765,N6745);
nand U2135 (N7800,N7787,N7769);
nand U2136 (N7803,N7788,N7771);
not U2137 (N7806,N7772);
nand U2138 (N7807,N7772,N6773);
not U2139 (N7808,N7775);
nand U2140 (N7809,N7775,N6777);
not U2141 (N7810,N7778);
nand U2142 (N7811,N7778,N6782);
nand U2143 (N7812,N7795,N7782);
nand U2144 (N7815,N6274,N7796);
nand U2145 (N7816,N6286,N7798);
nand U2146 (N7821,N6344,N7806);
nand U2147 (N7822,N6350,N7808);
nand U2148 (N7823,N6353,N7810);
nand U2149 (N7826,N7815,N7797);
nand U2150 (N7829,N7816,N7799);
not U2151 (N7832,N7800);
nand U2152 (N7833,N7800,N6752);
not U2153 (N7834,N7803);
nand U2154 (N7835,N7803,N6761);
nand U2155 (N7836,N7821,N7807);
nand U2156 (N7839,N7822,N7809);
nand U2157 (N7842,N7823,N7811);
not U2158 (N7845,N7812);
nand U2159 (N7846,N7812,N6790);
nand U2160 (N7851,N6298,N7832);
nand U2161 (N7852,N6316,N7834);
nand U2162 (N7859,N6364,N7845);
not U2163 (N7860,N7826);
nand U2164 (N7861,N7826,N6741);
not U2165 (N7862,N7829);
nand U2166 (N7863,N7829,N6746);
nand U2167 (N7864,N7851,N7833);
nand U2168 (N7867,N7852,N7835);
not U2169 (N7870,N7836);
nand U2170 (N7871,N7836,N5730);
not U2171 (N7872,N7839);
nand U2172 (N7873,N7839,N5732);
not U2173 (N7874,N7842);
nand U2174 (N7875,N7842,N6783);
nand U2175 (N7876,N7859,N7846);
nand U2176 (N7879,N6277,N7860);
nand U2177 (N7880,N6289,N7862);
nand U2178 (N7885,N5199,N7870);
nand U2179 (N7886,N5208,N7872);
nand U2180 (N7887,N6356,N7874);
nand U2181 (N7890,N7879,N7861);
nand U2182 (N7893,N7880,N7863);
not U2183 (N7896,N7864);
nand U2184 (N7897,N7864,N6753);
not U2185 (N7898,N7867);
nand U2186 (N7899,N7867,N6762);
nand U2187 (N7900,N7885,N7871);
nand U2188 (N7903,N7886,N7873);
nand U2189 (N7906,N7887,N7875);
not U2190 (N7909,N7876);
nand U2191 (N7910,N7876,N6791);
nand U2192 (N7917,N6301,N7896);
nand U2193 (N7918,N6319,N7898);
nand U2194 (N7923,N6367,N7909);
not U2195 (N7924,N7890);
nand U2196 (N7925,N7890,N6680);
not U2197 (N7926,N7893);
nand U2198 (N7927,N7893,N6681);
not U2199 (N7928,N7900);
nand U2200 (N7929,N7900,N5690);
not U2201 (N7930,N7903);
nand U2202 (N7931,N7903,N5691);
nand U2203 (N7932,N7917,N7897);
nand U2204 (N7935,N7918,N7899);
not U2205 (N7938,N7906);
nand U2206 (N7939,N7906,N6784);
nand U2207 (N7940,N7923,N7910);
nand U2208 (N7943,N6280,N7924);
nand U2209 (N7944,N6292,N7926);
nand U2210 (N7945,N5202,N7928);
nand U2211 (N7946,N5211,N7930);
nand U2212 (N7951,N6359,N7938);
nand U2213 (N7954,N7943,N7925);
nand U2214 (N7957,N7944,N7927);
nand U2215 (N7960,N7945,N7929);
nand U2216 (N7963,N7946,N7931);
not U2217 (N7966,N7932);
nand U2218 (N7967,N7932,N6754);
not U2219 (N7968,N7935);
nand U2220 (N7969,N7935,N6755);
nand U2221 (N7970,N7951,N7939);
not U2222 (N7973,N7940);
nand U2223 (N7974,N7940,N6785);
nand U2224 (N7984,N6304,N7966);
nand U2225 (N7985,N6322,N7968);
nand U2226 (N7987,N6370,N7973);
and U2227 (N7988,N7957,N6831,N1157);
and U2228 (N7989,N7954,N6415,N1157);
and U2229 (N7990,N7957,N7041,N566);
and U2230 (N7991,N7954,N7177,N566);
not U2231 (N7992,N7970);
nand U2232 (N7993,N7970,N6448);
and U2233 (N7994,N7963,N6857,N1219);
and U2234 (N7995,N7960,N6441,N1219);
and U2235 (N7996,N7963,N7065,N583);
and U2236 (N7997,N7960,N7182,N583);
nand U2237 (N7998,N7984,N7967);
nand U2238 (N8001,N7985,N7969);
nand U2239 (N8004,N7987,N7974);
nand U2240 (N8009,N6051,N7992);
or U2241 (N8013,N7988,N7989,N7990,N7991);
or U2242 (N8017,N7994,N7995,N7996,N7997);
not U2243 (N8020,N7998);
nand U2244 (N8021,N7998,N6682);
not U2245 (N8022,N8001);
nand U2246 (N8023,N8001,N6683);
nand U2247 (N8025,N8009,N7993);
not U2248 (N8026,N8004);
nand U2249 (N8027,N8004,N6449);
nand U2250 (N8031,N6307,N8020);
nand U2251 (N8032,N6310,N8022);
not U2252 (N8033,N8013);
nand U2253 (N8034,N6054,N8026);
and U2254 (N8035,N583,N8025);
not U2255 (N8036,N8017);
nand U2256 (N8037,N8031,N8021);
nand U2257 (N8038,N8032,N8023);
nand U2258 (N8039,N8034,N8027);
not U2259 (N8040,N8038);
and U2260 (N8041,N566,N8037);
not U2261 (N8042,N8039);
and U2262 (N8043,N8040,N1157);
and U2263 (N8044,N8042,N1219);
or U2264 (N8045,N8043,N8041);
or U2265 (N8048,N8044,N8035);
nand U2266 (N8055,N8045,N8033);
not U2267 (N8056,N8045);
nand U2268 (N8057,N8048,N8036);
not U2269 (N8058,N8048);
nand U2270 (N8059,N8013,N8056);
nand U2271 (N8060,N8017,N8058);
nand U2272 (N8061,N8055,N8059);
nand U2273 (N8064,N8057,N8060);
and U2274 (N8071,N8064,N1777,N3130);
and U2275 (N8072,N8061,N1761,N3108);
not U2276 (N8073,N8061);
not U2277 (N8074,N8064);
or U2278 (N8075,N7526,N8071,N3659,N2625);
or U2279 (N8076,N7636,N8072,N3661,N2627);
and U2280 (N8077,N8073,N1727);
and U2281 (N8078,N8074,N1727);
or U2282 (N8079,N7530,N8077);
or U2283 (N8082,N7479,N8078);
and U2284 (N8089,N8079,N3063);
and U2285 (N8090,N8082,N3063);
and U2286 (N8091,N8079,N3063);
and U2287 (N8092,N8082,N3063);
or U2288 (N8093,N8089,N3071);
or U2289 (N8096,N8090,N3072);
or U2290 (N8099,N8091,N3073);
or U2291 (N8102,N8092,N3074);
and U2292 (N8113,N8102,N2779,N2790);
and U2293 (N8114,N8099,N1327,N2790);
and U2294 (N8115,N8102,N2801,N2812);
and U2295 (N8116,N8099,N1351,N2812);
and U2296 (N8117,N8096,N2681,N2692);
and U2297 (N8118,N8093,N1185,N2692);
and U2298 (N8119,N8096,N2756,N2767);
and U2299 (N8120,N8093,N1247,N2767);
or U2300 (N8121,N8117,N8118,N3662,N2703);
or U2301 (N8122,N8119,N8120,N3663,N2778);
or U2302 (N8123,N8113,N8114,N3650,N2614);
or U2303 (N8124,N8115,N8116,N3658,N2622);
and U2304 (N8125,N8121,N2675);
and U2305 (N8126,N8122,N2750);
not U2306 (N8127,N8125);
not U2307 (N8128,N8126);
endmodule
