module c6288 (N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, N205, N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392, N409, N426, N443, N460, N477, N494, N511, N528, N545, N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, N5308, N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288);
input N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, N205, N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392, N409, N426, N443, N460, N477, N494, N511, N528;
output N545, N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, N5308, N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288;
wire N546, N549, N552, N555, N558, N561, N564, N567, N570, N573, N576, N579, N582, N585, N588, N591, N594, N597, N600, N603, N606, N609, N612, N615, N618, N621, N624, N627, N630, N633, N636, N639, N642, N645, N648, N651, N654, N657, N660, N663, N666, N669, N672, N675, N678, N681, N684, N687, N690, N693, N696, N699, N702, N705, N708, N711, N714, N717, N720, N723, N726, N729, N732, N735, N738, N741, N744, N747, N750, N753, N756, N759, N762, N765, N768, N771, N774, N777, N780, N783, N786, N789, N792, N795, N798, N801, N804, N807, N810, N813, N816, N819, N822, N825, N828, N831, N834, N837, N840, N843, N846, N849, N852, N855, N858, N861, N864, N867, N870, N873, N876, N879, N882, N885, N888, N891, N894, N897, N900, N903, N906, N909, N912, N915, N918, N921, N924, N927, N930, N933, N936, N939, N942, N945, N948, N951, N954, N957, N960, N963, N966, N969, N972, N975, N978, N981, N984, N987, N990, N993, N996, N999, N1002, N1005, N1008, N1011, N1014, N1017, N1020, N1023, N1026, N1029, N1032, N1035, N1038, N1041, N1044, N1047, N1050, N1053, N1056, N1059, N1062, N1065, N1068, N1071, N1074, N1077, N1080, N1083, N1086, N1089, N1092, N1095, N1098, N1101, N1104, N1107, N1110, N1113, N1116, N1119, N1122, N1125, N1128, N1131, N1134, N1137, N1140, N1143, N1146, N1149, N1152, N1155, N1158, N1161, N1164, N1167, N1170, N1173, N1176, N1179, N1182, N1185, N1188, N1191, N1194, N1197, N1200, N1203, N1206, N1209, N1212, N1215, N1218, N1221, N1224, N1227, N1230, N1233, N1236, N1239, N1242, N1245, N1248, N1251, N1254, N1257, N1260, N1263, N1266, N1269, N1272, N1275, N1278, N1281, N1284, N1287, N1290, N1293, N1296, N1299, N1302, N1305, N1308, N1311, N1315, N1319, N1323, N1327, N1331, N1335, N1339, N1343, N1347, N1351, N1355, N1359, N1363, N1367, N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394, N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1404, N1407, N1410, N1413, N1416, N1419, N1422, N1425, N1428, N1431, N1434, N1437, N1440, N1443, N1446, N1450, N1454, N1458, N1462, N1466, N1470, N1474, N1478, N1482, N1486, N1490, N1494, N1498, N1502, N1506, N1507, N1508, N1511, N1512, N1513, N1516, N1517, N1518, N1521, N1522, N1523, N1526, N1527, N1528, N1531, N1532, N1533, N1536, N1537, N1538, N1541, N1542, N1543, N1546, N1547, N1548, N1551, N1552, N1553, N1556, N1557, N1558, N1561, N1562, N1563, N1566, N1567, N1568, N1571, N1572, N1573, N1576, N1577, N1578, N1582, N1585, N1588, N1591, N1594, N1597, N1600, N1603, N1606, N1609, N1612, N1615, N1618, N1621, N1624, N1628, N1632, N1636, N1640, N1644, N1648, N1652, N1656, N1660, N1664, N1668, N1672, N1676, N1680, N1684, N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1692, N1693, N1694, N1695, N1696, N1697, N1698, N1699, N1700, N1701, N1702, N1703, N1704, N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712, N1713, N1714, N1717, N1720, N1723, N1726, N1729, N1732, N1735, N1738, N1741, N1744, N1747, N1750, N1753, N1756, N1759, N1763, N1767, N1771, N1775, N1779, N1783, N1787, N1791, N1795, N1799, N1803, N1807, N1811, N1815, N1819, N1820, N1821, N1824, N1825, N1826, N1829, N1830, N1831, N1834, N1835, N1836, N1839, N1840, N1841, N1844, N1845, N1846, N1849, N1850, N1851, N1854, N1855, N1856, N1859, N1860, N1861, N1864, N1865, N1866, N1869, N1870, N1871, N1874, N1875, N1876, N1879, N1880, N1881, N1884, N1885, N1886, N1889, N1890, N1891, N1894, N1897, N1902, N1905, N1908, N1911, N1914, N1917, N1920, N1923, N1926, N1929, N1932, N1935, N1938, N1941, N1945, N1946, N1947, N1951, N1955, N1959, N1963, N1967, N1971, N1975, N1979, N1983, N1987, N1991, N1995, N1999, N2000, N2001, N2004, N2005, N2006, N2007, N2008, N2009, N2010, N2011, N2012, N2013, N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024, N2025, N2026, N2027, N2028, N2029, N2030, N2033, N2037, N2040, N2043, N2046, N2049, N2052, N2055, N2058, N2061, N2064, N2067, N2070, N2073, N2076, N2080, N2081, N2082, N2085, N2089, N2093, N2097, N2101, N2105, N2109, N2113, N2117, N2121, N2125, N2129, N2133, N2137, N2138, N2139, N2142, N2145, N2149, N2150, N2151, N2154, N2155, N2156, N2159, N2160, N2161, N2164, N2165, N2166, N2169, N2170, N2171, N2174, N2175, N2176, N2179, N2180, N2181, N2184, N2185, N2186, N2189, N2190, N2191, N2194, N2195, N2196, N2199, N2200, N2201, N2204, N2205, N2206, N2209, N2210, N2211, N2214, N2217, N2221, N2222, N2224, N2227, N2230, N2233, N2236, N2239, N2242, N2245, N2248, N2251, N2254, N2257, N2260, N2264, N2265, N2266, N2269, N2273, N2277, N2281, N2285, N2289, N2293, N2297, N2301, N2305, N2309, N2313, N2317, N2318, N2319, N2322, N2326, N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338, N2339, N2340, N2341, N2342, N2343, N2344, N2345, N2346, N2347, N2348, N2349, N2350, N2353, N2357, N2358, N2359, N2362, N2365, N2368, N2371, N2374, N2377, N2380, N2383, N2386, N2389, N2392, N2395, N2398, N2402, N2403, N2404, N2407, N2410, N2414, N2418, N2422, N2426, N2430, N2434, N2438, N2442, N2446, N2450, N2454, N2458, N2462, N2463, N2464, N2467, N2470, N2474, N2475, N2476, N2477, N2478, N2481, N2482, N2483, N2486, N2487, N2488, N2491, N2492, N2493, N2496, N2497, N2498, N2501, N2502, N2503, N2506, N2507, N2508, N2511, N2512, N2513, N2516, N2517, N2518, N2521, N2522, N2523, N2526, N2527, N2528, N2531, N2532, N2533, N2536, N2539, N2543, N2544, N2545, N2549, N2552, N2555, N2558, N2561, N2564, N2567, N2570, N2573, N2576, N2579, N2582, N2586, N2587, N2588, N2591, N2595, N2599, N2603, N2607, N2611, N2615, N2619, N2623, N2627, N2631, N2635, N2639, N2640, N2641, N2644, N2648, N2649, N2650, N2653, N2654, N2655, N2656, N2657, N2658, N2659, N2660, N2661, N2662, N2663, N2664, N2665, N2666, N2667, N2668, N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2678, N2682, N2683, N2684, N2687, N2690, N2694, N2697, N2700, N2703, N2706, N2709, N2712, N2715, N2718, N2721, N2724, N2727, N2731, N2732, N2733, N2736, N2739, N2743, N2744, N2745, N2749, N2753, N2757, N2761, N2765, N2769, N2773, N2777, N2781, N2785, N2789, N2790, N2791, N2794, N2797, N2801, N2802, N2803, N2806, N2807, N2808, N2811, N2812, N2813, N2816, N2817, N2818, N2821, N2822, N2823, N2826, N2827, N2828, N2831, N2832, N2833, N2836, N2837, N2838, N2841, N2842, N2843, N2846, N2847, N2848, N2851, N2852, N2853, N2856, N2857, N2858, N2861, N2864, N2868, N2869, N2870, N2873, N2878, N2881, N2884, N2887, N2890, N2893, N2896, N2899, N2902, N2905, N2908, N2912, N2913, N2914, N2917, N2921, N2922, N2923, N2926, N2930, N2934, N2938, N2942, N2946, N2950, N2954, N2958, N2962, N2966, N2967, N2968, N2971, N2975, N2976, N2977, N2980, N2983, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005, N3006, N3007, N3010, N3014, N3015, N3016, N3019, N3022, N3026, N3027, N3028, N3031, N3034, N3037, N3040, N3043, N3046, N3049, N3052, N3055, N3058, N3062, N3063, N3064, N3067, N3070, N3074, N3075, N3076, N3079, N3083, N3087, N3091, N3095, N3099, N3103, N3107, N3111, N3115, N3119, N3120, N3121, N3124, N3127, N3131, N3132, N3133, N3136, N3140, N3141, N3142, N3145, N3146, N3147, N3150, N3151, N3152, N3155, N3156, N3157, N3160, N3161, N3162, N3165, N3166, N3167, N3170, N3171, N3172, N3175, N3176, N3177, N3180, N3181, N3182, N3185, N3186, N3187, N3190, N3193, N3197, N3198, N3199, N3202, N3206, N3207, N3208, N3212, N3215, N3218, N3221, N3224, N3227, N3230, N3233, N3236, N3239, N3243, N3244, N3245, N3248, N3252, N3253, N3254, N3257, N3260, N3264, N3268, N3272, N3276, N3280, N3284, N3288, N3292, N3296, N3300, N3301, N3302, N3305, N3309, N3310, N3311, N3314, N3317, N3321, N3322, N3323, N3324, N3325, N3326, N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334, N3335, N3336, N3337, N3338, N3339, N3340, N3341, N3344, N3348, N3349, N3350, N3353, N3356, N3360, N3361, N3362, N3365, N3368, N3371, N3374, N3377, N3380, N3383, N3386, N3389, N3392, N3396, N3397, N3398, N3401, N3404, N3408, N3409, N3410, N3413, N3417, N3421, N3425, N3429, N3433, N3437, N3441, N3445, N3449, N3453, N3454, N3455, N3458, N3461, N3465, N3466, N3467, N3470, N3474, N3475, N3476, N3479, N3480, N3481, N3484, N3485, N3486, N3489, N3490, N3491, N3494, N3495, N3496, N3499, N3500, N3501, N3504, N3505, N3506, N3509, N3510, N3511, N3514, N3515, N3516, N3519, N3520, N3521, N3524, N3527, N3531, N3532, N3533, N3536, N3540, N3541, N3542, N3545, N3548, N3553, N3556, N3559, N3562, N3565, N3568, N3571, N3574, N3577, N3581, N3582, N3583, N3586, N3590, N3591, N3592, N3595, N3598, N3602, N3603, N3604, N3608, N3612, N3616, N3620, N3624, N3628, N3632, N3636, N3637, N3638, N3641, N3645, N3646, N3647, N3650, N3653, N3657, N3658, N3659, N3662, N3663, N3664, N3665, N3666, N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676, N3677, N3678, N3681, N3685, N3686, N3687, N3690, N3693, N3697, N3698, N3699, N3702, N3706, N3709, N3712, N3715, N3718, N3721, N3724, N3727, N3730, N3734, N3735, N3736, N3739, N3742, N3746, N3747, N3748, N3751, N3755, N3756, N3757, N3760, N3764, N3768, N3772, N3776, N3780, N3784, N3788, N3792, N3793, N3794, N3797, N3800, N3804, N3805, N3806, N3809, N3813, N3814, N3815, N3818, N3821, N3825, N3826, N3827, N3830, N3831, N3832, N3835, N3836, N3837, N3840, N3841, N3842, N3845, N3846, N3847, N3850, N3851, N3852, N3855, N3856, N3857, N3860, N3861, N3862, N3865, N3868, N3872, N3873, N3874, N3877, N3881, N3882, N3883, N3886, N3889, N3893, N3894, N3896, N3899, N3902, N3905, N3908, N3911, N3914, N3917, N3921, N3922, N3923, N3926, N3930, N3931, N3932, N3935, N3938, N3942, N3943, N3944, N3947, N3951, N3955, N3959, N3963, N3967, N3971, N3975, N3976, N3977, N3980, N3984, N3985, N3986, N3989, N3992, N3996, N3997, N3998, N4001, N4005, N4006, N4007, N4008, N4009, N4010, N4011, N4012, N4013, N4014, N4015, N4016, N4017, N4018, N4019, N4022, N4026, N4027, N4028, N4031, N4034, N4038, N4039, N4040, N4043, N4047, N4048, N4049, N4052, N4055, N4058, N4061, N4064, N4067, N4070, N4073, N4077, N4078, N4079, N4082, N4085, N4089, N4090, N4091, N4094, N4098, N4099, N4100, N4103, N4106, N4110, N4114, N4118, N4122, N4126, N4130, N4134, N4138, N4139, N4140, N4143, N4146, N4150, N4151, N4152, N4155, N4159, N4160, N4161, N4164, N4167, N4171, N4172, N4173, N4174, N4175, N4178, N4179, N4180, N4183, N4184, N4185, N4188, N4189, N4190, N4193, N4194, N4195, N4198, N4199, N4200, N4203, N4204, N4205, N4208, N4211, N4215, N4216, N4217, N4220, N4224, N4225, N4226, N4229, N4232, N4236, N4237, N4238, N4242, N4245, N4248, N4251, N4254, N4257, N4260, N4264, N4265, N4266, N4269, N4273, N4274, N4275, N4278, N4281, N4285, N4286, N4287, N4290, N4294, N4298, N4302, N4306, N4310, N4314, N4318, N4319, N4320, N4323, N4327, N4328, N4329, N4332, N4335, N4339, N4340, N4341, N4344, N4348, N4349, N4350, N4353, N4354, N4355, N4356, N4357, N4358, N4359, N4360, N4361, N4362, N4363, N4364, N4365, N4368, N4372, N4373, N4374, N4377, N4380, N4384, N4385, N4386, N4389, N4393, N4394, N4395, N4398, N4401, N4405, N4408, N4411, N4414, N4417, N4420, N4423, N4427, N4428, N4429, N4432, N4435, N4439, N4440, N4441, N4444, N4448, N4449, N4450, N4453, N4456, N4460, N4461, N4462, N4466, N4470, N4474, N4478, N4482, N4486, N4487, N4488, N4491, N4494, N4498, N4499, N4500, N4503, N4507, N4508, N4509, N4512, N4515, N4519, N4520, N4521, N4524, N4525, N4526, N4529, N4530, N4531, N4534, N4535, N4536, N4539, N4540, N4541, N4544, N4545, N4546, N4549, N4550, N4551, N4554, N4557, N4561, N4562, N4563, N4566, N4570, N4571, N4572, N4575, N4578, N4582, N4583, N4584, N4587, N4592, N4595, N4598, N4601, N4604, N4607, N4611, N4612, N4613, N4616, N4620, N4621, N4622, N4625, N4628, N4632, N4633, N4634, N4637, N4641, N4642, N4643, N4646, N4650, N4654, N4658, N4662, N4666, N4667, N4668, N4671, N4675, N4676, N4677, N4680, N4683, N4687, N4688, N4689, N4692, N4696, N4697, N4698, N4701, N4704, N4708, N4709, N4710, N4711, N4712, N4713, N4714, N4715, N4716, N4717, N4718, N4721, N4725, N4726, N4727, N4730, N4733, N4737, N4738, N4739, N4742, N4746, N4747, N4748, N4751, N4754, N4758, N4759, N4760, N4763, N4766, N4769, N4772, N4775, N4779, N4780, N4781, N4784, N4787, N4791, N4792, N4793, N4796, N4800, N4801, N4802, N4805, N4808, N4812, N4813, N4814, N4817, N4821, N4825, N4829, N4833, N4837, N4838, N4839, N4842, N4845, N4849, N4850, N4851, N4854, N4858, N4859, N4860, N4863, N4866, N4870, N4871, N4872, N4875, N4879, N4880, N4881, N4884, N4885, N4886, N4889, N4890, N4891, N4894, N4895, N4896, N4899, N4900, N4901, N4904, N4907, N4911, N4912, N4913, N4916, N4920, N4921, N4922, N4925, N4928, N4932, N4933, N4934, N4937, N4941, N4942, N4943, N4947, N4950, N4953, N4956, N4959, N4963, N4964, N4965, N4968, N4972, N4973, N4974, N4977, N4980, N4984, N4985, N4986, N4989, N4993, N4994, N4995, N4998, N5001, N5005, N5009, N5013, N5017, N5021, N5022, N5023, N5026, N5030, N5031, N5032, N5035, N5038, N5042, N5043, N5044, N5047, N5051, N5052, N5053, N5056, N5059, N5063, N5064, N5065, N5066, N5067, N5068, N5069, N5070, N5071, N5072, N5073, N5076, N5080, N5081, N5082, N5085, N5088, N5092, N5093, N5094, N5097, N5101, N5102, N5103, N5106, N5109, N5113, N5114, N5115, N5118, N5121, N5124, N5127, N5130, N5134, N5135, N5136, N5139, N5142, N5146, N5147, N5148, N5151, N5155, N5156, N5157, N5160, N5163, N5167, N5168, N5169, N5172, N5176, N5180, N5184, N5188, N5192, N5193, N5194, N5197, N5200, N5204, N5205, N5206, N5209, N5213, N5214, N5215, N5218, N5221, N5225, N5226, N5227, N5230, N5234, N5235, N5236, N5239, N5240, N5241, N5244, N5245, N5246, N5249, N5250, N5251, N5254, N5255, N5256, N5259, N5262, N5266, N5267, N5268, N5271, N5275, N5276, N5277, N5280, N5283, N5287, N5288, N5289, N5292, N5296, N5297, N5298, N5301, N5304, N5309, N5312, N5315, N5318, N5322, N5323, N5324, N5327, N5331, N5332, N5333, N5336, N5339, N5343, N5344, N5345, N5348, N5352, N5353, N5354, N5357, N5360, N5364, N5365, N5366, N5370, N5374, N5378, N5379, N5380, N5383, N5387, N5388, N5389, N5392, N5395, N5399, N5400, N5401, N5404, N5408, N5409, N5410, N5413, N5416, N5420, N5421, N5422, N5425, N5426, N5427, N5428, N5429, N5430, N5431, N5434, N5438, N5439, N5440, N5443, N5446, N5450, N5451, N5452, N5455, N5459, N5460, N5461, N5464, N5467, N5471, N5472, N5473, N5476, N5480, N5483, N5486, N5489, N5493, N5494, N5495, N5498, N5501, N5505, N5506, N5507, N5510, N5514, N5515, N5516, N5519, N5522, N5526, N5527, N5528, N5531, N5535, N5536, N5537, N5540, N5544, N5548, N5552, N5553, N5554, N5557, N5560, N5564, N5565, N5566, N5569, N5573, N5574, N5575, N5578, N5581, N5585, N5586, N5587, N5590, N5594, N5595, N5596, N5599, N5602, N5606, N5607, N5608, N5611, N5612, N5613, N5616, N5617, N5618, N5621, N5624, N5628, N5629, N5630, N5633, N5637, N5638, N5639, N5642, N5645, N5649, N5650, N5651, N5654, N5658, N5659, N5660, N5663, N5666, N5670, N5671, N5673, N5676, N5679, N5683, N5684, N5685, N5688, N5692, N5693, N5694, N5697, N5700, N5704, N5705, N5706, N5709, N5713, N5714, N5715, N5718, N5721, N5725, N5726, N5727, N5730, N5734, N5738, N5739, N5740, N5743, N5747, N5748, N5749, N5752, N5755, N5759, N5760, N5761, N5764, N5768, N5769, N5770, N5773, N5776, N5780, N5781, N5782, N5785, N5786, N5787, N5788, N5789, N5792, N5796, N5797, N5798, N5801, N5804, N5808, N5809, N5810, N5813, N5817, N5818, N5819, N5822, N5825, N5829, N5830, N5831, N5834, N5837, N5840, N5844, N5845, N5846, N5849, N5852, N5856, N5857, N5858, N5861, N5865, N5866, N5867, N5870, N5873, N5877, N5878, N5879, N5882, N5886, N5890, N5891, N5892, N5895, N5898, N5902, N5903, N5904, N5907, N5911, N5912, N5913, N5916, N5919, N5923, N5924, N5925, N5928, N5929, N5930, N5933, N5934, N5935, N5938, N5941, N5945, N5946, N5947, N5950, N5954, N5955, N5956, N5959, N5962, N5966, N5967, N5968, N5972, N5975, N5979, N5980, N5981, N5984, N5988, N5989, N5990, N5993, N5996, N6000, N6001, N6002, N6005, N6009, N6010, N6011, N6014, N6018, N6019, N6020, N6023, N6026, N6030, N6031, N6032, N6035, N6036, N6037, N6040, N6044, N6045, N6046, N6049, N6052, N6056, N6057, N6058, N6061, N6064, N6068, N6069, N6070, N6073, N6076, N6080, N6081, N6082, N6085, N6089, N6090, N6091, N6094, N6097, N6101, N6102, N6103, N6106, N6107, N6108, N6111, N6114, N6118, N6119, N6120, N6124, N6128, N6129, N6130, N6133, N6134, N6135, N6138, N6141, N6145, N6146, N6147, N6151, N6155, N6156, N6157, N6161, N6165, N6166, N6167, N6171, N6175, N6176, N6177, N6181, N6185, N6186, N6187, N6191, N6195, N6196, N6197, N6201, N6205, N6206, N6207, N6211, N6215, N6216, N6217, N6221, N6225, N6226, N6227, N6231, N6235, N6236, N6237, N6241, N6245, N6246, N6247, N6251, N6255, N6256, N6257, N6261, N6265, N6266, N6267, N6271, N6275, N6276, N6277, N6281, N6285, N6286;

and U1 (N545,N1,N273);
and U2 (N546,N1,N290);
and U3 (N549,N1,N307);
and U4 (N552,N1,N324);
and U5 (N555,N1,N341);
and U6 (N558,N1,N358);
and U7 (N561,N1,N375);
and U8 (N564,N1,N392);
and U9 (N567,N1,N409);
and U10 (N570,N1,N426);
and U11 (N573,N1,N443);
and U12 (N576,N1,N460);
and U13 (N579,N1,N477);
and U14 (N582,N1,N494);
and U15 (N585,N1,N511);
and U16 (N588,N1,N528);
and U17 (N591,N18,N273);
and U18 (N594,N18,N290);
and U19 (N597,N18,N307);
and U20 (N600,N18,N324);
and U21 (N603,N18,N341);
and U22 (N606,N18,N358);
and U23 (N609,N18,N375);
and U24 (N612,N18,N392);
and U25 (N615,N18,N409);
and U26 (N618,N18,N426);
and U27 (N621,N18,N443);
and U28 (N624,N18,N460);
and U29 (N627,N18,N477);
and U30 (N630,N18,N494);
and U31 (N633,N18,N511);
and U32 (N636,N18,N528);
and U33 (N639,N35,N273);
and U34 (N642,N35,N290);
and U35 (N645,N35,N307);
and U36 (N648,N35,N324);
and U37 (N651,N35,N341);
and U38 (N654,N35,N358);
and U39 (N657,N35,N375);
and U40 (N660,N35,N392);
and U41 (N663,N35,N409);
and U42 (N666,N35,N426);
and U43 (N669,N35,N443);
and U44 (N672,N35,N460);
and U45 (N675,N35,N477);
and U46 (N678,N35,N494);
and U47 (N681,N35,N511);
and U48 (N684,N35,N528);
and U49 (N687,N52,N273);
and U50 (N690,N52,N290);
and U51 (N693,N52,N307);
and U52 (N696,N52,N324);
and U53 (N699,N52,N341);
and U54 (N702,N52,N358);
and U55 (N705,N52,N375);
and U56 (N708,N52,N392);
and U57 (N711,N52,N409);
and U58 (N714,N52,N426);
and U59 (N717,N52,N443);
and U60 (N720,N52,N460);
and U61 (N723,N52,N477);
and U62 (N726,N52,N494);
and U63 (N729,N52,N511);
and U64 (N732,N52,N528);
and U65 (N735,N69,N273);
and U66 (N738,N69,N290);
and U67 (N741,N69,N307);
and U68 (N744,N69,N324);
and U69 (N747,N69,N341);
and U70 (N750,N69,N358);
and U71 (N753,N69,N375);
and U72 (N756,N69,N392);
and U73 (N759,N69,N409);
and U74 (N762,N69,N426);
and U75 (N765,N69,N443);
and U76 (N768,N69,N460);
and U77 (N771,N69,N477);
and U78 (N774,N69,N494);
and U79 (N777,N69,N511);
and U80 (N780,N69,N528);
and U81 (N783,N86,N273);
and U82 (N786,N86,N290);
and U83 (N789,N86,N307);
and U84 (N792,N86,N324);
and U85 (N795,N86,N341);
and U86 (N798,N86,N358);
and U87 (N801,N86,N375);
and U88 (N804,N86,N392);
and U89 (N807,N86,N409);
and U90 (N810,N86,N426);
and U91 (N813,N86,N443);
and U92 (N816,N86,N460);
and U93 (N819,N86,N477);
and U94 (N822,N86,N494);
and U95 (N825,N86,N511);
and U96 (N828,N86,N528);
and U97 (N831,N103,N273);
and U98 (N834,N103,N290);
and U99 (N837,N103,N307);
and U100 (N840,N103,N324);
and U101 (N843,N103,N341);
and U102 (N846,N103,N358);
and U103 (N849,N103,N375);
and U104 (N852,N103,N392);
and U105 (N855,N103,N409);
and U106 (N858,N103,N426);
and U107 (N861,N103,N443);
and U108 (N864,N103,N460);
and U109 (N867,N103,N477);
and U110 (N870,N103,N494);
and U111 (N873,N103,N511);
and U112 (N876,N103,N528);
and U113 (N879,N120,N273);
and U114 (N882,N120,N290);
and U115 (N885,N120,N307);
and U116 (N888,N120,N324);
and U117 (N891,N120,N341);
and U118 (N894,N120,N358);
and U119 (N897,N120,N375);
and U120 (N900,N120,N392);
and U121 (N903,N120,N409);
and U122 (N906,N120,N426);
and U123 (N909,N120,N443);
and U124 (N912,N120,N460);
and U125 (N915,N120,N477);
and U126 (N918,N120,N494);
and U127 (N921,N120,N511);
and U128 (N924,N120,N528);
and U129 (N927,N137,N273);
and U130 (N930,N137,N290);
and U131 (N933,N137,N307);
and U132 (N936,N137,N324);
and U133 (N939,N137,N341);
and U134 (N942,N137,N358);
and U135 (N945,N137,N375);
and U136 (N948,N137,N392);
and U137 (N951,N137,N409);
and U138 (N954,N137,N426);
and U139 (N957,N137,N443);
and U140 (N960,N137,N460);
and U141 (N963,N137,N477);
and U142 (N966,N137,N494);
and U143 (N969,N137,N511);
and U144 (N972,N137,N528);
and U145 (N975,N154,N273);
and U146 (N978,N154,N290);
and U147 (N981,N154,N307);
and U148 (N984,N154,N324);
and U149 (N987,N154,N341);
and U150 (N990,N154,N358);
and U151 (N993,N154,N375);
and U152 (N996,N154,N392);
and U153 (N999,N154,N409);
and U154 (N1002,N154,N426);
and U155 (N1005,N154,N443);
and U156 (N1008,N154,N460);
and U157 (N1011,N154,N477);
and U158 (N1014,N154,N494);
and U159 (N1017,N154,N511);
and U160 (N1020,N154,N528);
and U161 (N1023,N171,N273);
and U162 (N1026,N171,N290);
and U163 (N1029,N171,N307);
and U164 (N1032,N171,N324);
and U165 (N1035,N171,N341);
and U166 (N1038,N171,N358);
and U167 (N1041,N171,N375);
and U168 (N1044,N171,N392);
and U169 (N1047,N171,N409);
and U170 (N1050,N171,N426);
and U171 (N1053,N171,N443);
and U172 (N1056,N171,N460);
and U173 (N1059,N171,N477);
and U174 (N1062,N171,N494);
and U175 (N1065,N171,N511);
and U176 (N1068,N171,N528);
and U177 (N1071,N188,N273);
and U178 (N1074,N188,N290);
and U179 (N1077,N188,N307);
and U180 (N1080,N188,N324);
and U181 (N1083,N188,N341);
and U182 (N1086,N188,N358);
and U183 (N1089,N188,N375);
and U184 (N1092,N188,N392);
and U185 (N1095,N188,N409);
and U186 (N1098,N188,N426);
and U187 (N1101,N188,N443);
and U188 (N1104,N188,N460);
and U189 (N1107,N188,N477);
and U190 (N1110,N188,N494);
and U191 (N1113,N188,N511);
and U192 (N1116,N188,N528);
and U193 (N1119,N205,N273);
and U194 (N1122,N205,N290);
and U195 (N1125,N205,N307);
and U196 (N1128,N205,N324);
and U197 (N1131,N205,N341);
and U198 (N1134,N205,N358);
and U199 (N1137,N205,N375);
and U200 (N1140,N205,N392);
and U201 (N1143,N205,N409);
and U202 (N1146,N205,N426);
and U203 (N1149,N205,N443);
and U204 (N1152,N205,N460);
and U205 (N1155,N205,N477);
and U206 (N1158,N205,N494);
and U207 (N1161,N205,N511);
and U208 (N1164,N205,N528);
and U209 (N1167,N222,N273);
and U210 (N1170,N222,N290);
and U211 (N1173,N222,N307);
and U212 (N1176,N222,N324);
and U213 (N1179,N222,N341);
and U214 (N1182,N222,N358);
and U215 (N1185,N222,N375);
and U216 (N1188,N222,N392);
and U217 (N1191,N222,N409);
and U218 (N1194,N222,N426);
and U219 (N1197,N222,N443);
and U220 (N1200,N222,N460);
and U221 (N1203,N222,N477);
and U222 (N1206,N222,N494);
and U223 (N1209,N222,N511);
and U224 (N1212,N222,N528);
and U225 (N1215,N239,N273);
and U226 (N1218,N239,N290);
and U227 (N1221,N239,N307);
and U228 (N1224,N239,N324);
and U229 (N1227,N239,N341);
and U230 (N1230,N239,N358);
and U231 (N1233,N239,N375);
and U232 (N1236,N239,N392);
and U233 (N1239,N239,N409);
and U234 (N1242,N239,N426);
and U235 (N1245,N239,N443);
and U236 (N1248,N239,N460);
and U237 (N1251,N239,N477);
and U238 (N1254,N239,N494);
and U239 (N1257,N239,N511);
and U240 (N1260,N239,N528);
and U241 (N1263,N256,N273);
and U242 (N1266,N256,N290);
and U243 (N1269,N256,N307);
and U244 (N1272,N256,N324);
and U245 (N1275,N256,N341);
and U246 (N1278,N256,N358);
and U247 (N1281,N256,N375);
and U248 (N1284,N256,N392);
and U249 (N1287,N256,N409);
and U250 (N1290,N256,N426);
and U251 (N1293,N256,N443);
and U252 (N1296,N256,N460);
and U253 (N1299,N256,N477);
and U254 (N1302,N256,N494);
and U255 (N1305,N256,N511);
and U256 (N1308,N256,N528);
not U257 (N1311,N591);
not U258 (N1315,N639);
not U259 (N1319,N687);
not U260 (N1323,N735);
not U261 (N1327,N783);
not U262 (N1331,N831);
not U263 (N1335,N879);
not U264 (N1339,N927);
not U265 (N1343,N975);
not U266 (N1347,N1023);
not U267 (N1351,N1071);
not U268 (N1355,N1119);
not U269 (N1359,N1167);
not U270 (N1363,N1215);
not U271 (N1367,N1263);
nor U272 (N1371,N591,N1311);
not U273 (N1372,N1311);
nor U274 (N1373,N639,N1315);
not U275 (N1374,N1315);
nor U276 (N1375,N687,N1319);
not U277 (N1376,N1319);
nor U278 (N1377,N735,N1323);
not U279 (N1378,N1323);
nor U280 (N1379,N783,N1327);
not U281 (N1380,N1327);
nor U282 (N1381,N831,N1331);
not U283 (N1382,N1331);
nor U284 (N1383,N879,N1335);
not U285 (N1384,N1335);
nor U286 (N1385,N927,N1339);
not U287 (N1386,N1339);
nor U288 (N1387,N975,N1343);
not U289 (N1388,N1343);
nor U290 (N1389,N1023,N1347);
not U291 (N1390,N1347);
nor U292 (N1391,N1071,N1351);
not U293 (N1392,N1351);
nor U294 (N1393,N1119,N1355);
not U295 (N1394,N1355);
nor U296 (N1395,N1167,N1359);
not U297 (N1396,N1359);
nor U298 (N1397,N1215,N1363);
not U299 (N1398,N1363);
nor U300 (N1399,N1263,N1367);
not U301 (N1400,N1367);
nor U302 (N1401,N1371,N1372);
nor U303 (N1404,N1373,N1374);
nor U304 (N1407,N1375,N1376);
nor U305 (N1410,N1377,N1378);
nor U306 (N1413,N1379,N1380);
nor U307 (N1416,N1381,N1382);
nor U308 (N1419,N1383,N1384);
nor U309 (N1422,N1385,N1386);
nor U310 (N1425,N1387,N1388);
nor U311 (N1428,N1389,N1390);
nor U312 (N1431,N1391,N1392);
nor U313 (N1434,N1393,N1394);
nor U314 (N1437,N1395,N1396);
nor U315 (N1440,N1397,N1398);
nor U316 (N1443,N1399,N1400);
nor U317 (N1446,N1401,N546);
nor U318 (N1450,N1404,N594);
nor U319 (N1454,N1407,N642);
nor U320 (N1458,N1410,N690);
nor U321 (N1462,N1413,N738);
nor U322 (N1466,N1416,N786);
nor U323 (N1470,N1419,N834);
nor U324 (N1474,N1422,N882);
nor U325 (N1478,N1425,N930);
nor U326 (N1482,N1428,N978);
nor U327 (N1486,N1431,N1026);
nor U328 (N1490,N1434,N1074);
nor U329 (N1494,N1437,N1122);
nor U330 (N1498,N1440,N1170);
nor U331 (N1502,N1443,N1218);
nor U332 (N1506,N1401,N1446);
nor U333 (N1507,N1446,N546);
nor U334 (N1508,N1311,N1446);
nor U335 (N1511,N1404,N1450);
nor U336 (N1512,N1450,N594);
nor U337 (N1513,N1315,N1450);
nor U338 (N1516,N1407,N1454);
nor U339 (N1517,N1454,N642);
nor U340 (N1518,N1319,N1454);
nor U341 (N1521,N1410,N1458);
nor U342 (N1522,N1458,N690);
nor U343 (N1523,N1323,N1458);
nor U344 (N1526,N1413,N1462);
nor U345 (N1527,N1462,N738);
nor U346 (N1528,N1327,N1462);
nor U347 (N1531,N1416,N1466);
nor U348 (N1532,N1466,N786);
nor U349 (N1533,N1331,N1466);
nor U350 (N1536,N1419,N1470);
nor U351 (N1537,N1470,N834);
nor U352 (N1538,N1335,N1470);
nor U353 (N1541,N1422,N1474);
nor U354 (N1542,N1474,N882);
nor U355 (N1543,N1339,N1474);
nor U356 (N1546,N1425,N1478);
nor U357 (N1547,N1478,N930);
nor U358 (N1548,N1343,N1478);
nor U359 (N1551,N1428,N1482);
nor U360 (N1552,N1482,N978);
nor U361 (N1553,N1347,N1482);
nor U362 (N1556,N1431,N1486);
nor U363 (N1557,N1486,N1026);
nor U364 (N1558,N1351,N1486);
nor U365 (N1561,N1434,N1490);
nor U366 (N1562,N1490,N1074);
nor U367 (N1563,N1355,N1490);
nor U368 (N1566,N1437,N1494);
nor U369 (N1567,N1494,N1122);
nor U370 (N1568,N1359,N1494);
nor U371 (N1571,N1440,N1498);
nor U372 (N1572,N1498,N1170);
nor U373 (N1573,N1363,N1498);
nor U374 (N1576,N1443,N1502);
nor U375 (N1577,N1502,N1218);
nor U376 (N1578,N1367,N1502);
nor U377 (N1581,N1506,N1507);
nor U378 (N1582,N1511,N1512);
nor U379 (N1585,N1516,N1517);
nor U380 (N1588,N1521,N1522);
nor U381 (N1591,N1526,N1527);
nor U382 (N1594,N1531,N1532);
nor U383 (N1597,N1536,N1537);
nor U384 (N1600,N1541,N1542);
nor U385 (N1603,N1546,N1547);
nor U386 (N1606,N1551,N1552);
nor U387 (N1609,N1556,N1557);
nor U388 (N1612,N1561,N1562);
nor U389 (N1615,N1566,N1567);
nor U390 (N1618,N1571,N1572);
nor U391 (N1621,N1576,N1577);
nor U392 (N1624,N1266,N1578);
nor U393 (N1628,N1582,N1508);
nor U394 (N1632,N1585,N1513);
nor U395 (N1636,N1588,N1518);
nor U396 (N1640,N1591,N1523);
nor U397 (N1644,N1594,N1528);
nor U398 (N1648,N1597,N1533);
nor U399 (N1652,N1600,N1538);
nor U400 (N1656,N1603,N1543);
nor U401 (N1660,N1606,N1548);
nor U402 (N1664,N1609,N1553);
nor U403 (N1668,N1612,N1558);
nor U404 (N1672,N1615,N1563);
nor U405 (N1676,N1618,N1568);
nor U406 (N1680,N1621,N1573);
nor U407 (N1684,N1266,N1624);
nor U408 (N1685,N1624,N1578);
nor U409 (N1686,N1582,N1628);
nor U410 (N1687,N1628,N1508);
nor U411 (N1688,N1585,N1632);
nor U412 (N1689,N1632,N1513);
nor U413 (N1690,N1588,N1636);
nor U414 (N1691,N1636,N1518);
nor U415 (N1692,N1591,N1640);
nor U416 (N1693,N1640,N1523);
nor U417 (N1694,N1594,N1644);
nor U418 (N1695,N1644,N1528);
nor U419 (N1696,N1597,N1648);
nor U420 (N1697,N1648,N1533);
nor U421 (N1698,N1600,N1652);
nor U422 (N1699,N1652,N1538);
nor U423 (N1700,N1603,N1656);
nor U424 (N1701,N1656,N1543);
nor U425 (N1702,N1606,N1660);
nor U426 (N1703,N1660,N1548);
nor U427 (N1704,N1609,N1664);
nor U428 (N1705,N1664,N1553);
nor U429 (N1706,N1612,N1668);
nor U430 (N1707,N1668,N1558);
nor U431 (N1708,N1615,N1672);
nor U432 (N1709,N1672,N1563);
nor U433 (N1710,N1618,N1676);
nor U434 (N1711,N1676,N1568);
nor U435 (N1712,N1621,N1680);
nor U436 (N1713,N1680,N1573);
nor U437 (N1714,N1684,N1685);
nor U438 (N1717,N1686,N1687);
nor U439 (N1720,N1688,N1689);
nor U440 (N1723,N1690,N1691);
nor U441 (N1726,N1692,N1693);
nor U442 (N1729,N1694,N1695);
nor U443 (N1732,N1696,N1697);
nor U444 (N1735,N1698,N1699);
nor U445 (N1738,N1700,N1701);
nor U446 (N1741,N1702,N1703);
nor U447 (N1744,N1704,N1705);
nor U448 (N1747,N1706,N1707);
nor U449 (N1750,N1708,N1709);
nor U450 (N1753,N1710,N1711);
nor U451 (N1756,N1712,N1713);
nor U452 (N1759,N1714,N1221);
nor U453 (N1763,N1717,N549);
nor U454 (N1767,N1720,N597);
nor U455 (N1771,N1723,N645);
nor U456 (N1775,N1726,N693);
nor U457 (N1779,N1729,N741);
nor U458 (N1783,N1732,N789);
nor U459 (N1787,N1735,N837);
nor U460 (N1791,N1738,N885);
nor U461 (N1795,N1741,N933);
nor U462 (N1799,N1744,N981);
nor U463 (N1803,N1747,N1029);
nor U464 (N1807,N1750,N1077);
nor U465 (N1811,N1753,N1125);
nor U466 (N1815,N1756,N1173);
nor U467 (N1819,N1714,N1759);
nor U468 (N1820,N1759,N1221);
nor U469 (N1821,N1624,N1759);
nor U470 (N1824,N1717,N1763);
nor U471 (N1825,N1763,N549);
nor U472 (N1826,N1628,N1763);
nor U473 (N1829,N1720,N1767);
nor U474 (N1830,N1767,N597);
nor U475 (N1831,N1632,N1767);
nor U476 (N1834,N1723,N1771);
nor U477 (N1835,N1771,N645);
nor U478 (N1836,N1636,N1771);
nor U479 (N1839,N1726,N1775);
nor U480 (N1840,N1775,N693);
nor U481 (N1841,N1640,N1775);
nor U482 (N1844,N1729,N1779);
nor U483 (N1845,N1779,N741);
nor U484 (N1846,N1644,N1779);
nor U485 (N1849,N1732,N1783);
nor U486 (N1850,N1783,N789);
nor U487 (N1851,N1648,N1783);
nor U488 (N1854,N1735,N1787);
nor U489 (N1855,N1787,N837);
nor U490 (N1856,N1652,N1787);
nor U491 (N1859,N1738,N1791);
nor U492 (N1860,N1791,N885);
nor U493 (N1861,N1656,N1791);
nor U494 (N1864,N1741,N1795);
nor U495 (N1865,N1795,N933);
nor U496 (N1866,N1660,N1795);
nor U497 (N1869,N1744,N1799);
nor U498 (N1870,N1799,N981);
nor U499 (N1871,N1664,N1799);
nor U500 (N1874,N1747,N1803);
nor U501 (N1875,N1803,N1029);
nor U502 (N1876,N1668,N1803);
nor U503 (N1879,N1750,N1807);
nor U504 (N1880,N1807,N1077);
nor U505 (N1881,N1672,N1807);
nor U506 (N1884,N1753,N1811);
nor U507 (N1885,N1811,N1125);
nor U508 (N1886,N1676,N1811);
nor U509 (N1889,N1756,N1815);
nor U510 (N1890,N1815,N1173);
nor U511 (N1891,N1680,N1815);
nor U512 (N1894,N1819,N1820);
nor U513 (N1897,N1269,N1821);
nor U514 (N1901,N1824,N1825);
nor U515 (N1902,N1829,N1830);
nor U516 (N1905,N1834,N1835);
nor U517 (N1908,N1839,N1840);
nor U518 (N1911,N1844,N1845);
nor U519 (N1914,N1849,N1850);
nor U520 (N1917,N1854,N1855);
nor U521 (N1920,N1859,N1860);
nor U522 (N1923,N1864,N1865);
nor U523 (N1926,N1869,N1870);
nor U524 (N1929,N1874,N1875);
nor U525 (N1932,N1879,N1880);
nor U526 (N1935,N1884,N1885);
nor U527 (N1938,N1889,N1890);
nor U528 (N1941,N1894,N1891);
nor U529 (N1945,N1269,N1897);
nor U530 (N1946,N1897,N1821);
nor U531 (N1947,N1902,N1826);
nor U532 (N1951,N1905,N1831);
nor U533 (N1955,N1908,N1836);
nor U534 (N1959,N1911,N1841);
nor U535 (N1963,N1914,N1846);
nor U536 (N1967,N1917,N1851);
nor U537 (N1971,N1920,N1856);
nor U538 (N1975,N1923,N1861);
nor U539 (N1979,N1926,N1866);
nor U540 (N1983,N1929,N1871);
nor U541 (N1987,N1932,N1876);
nor U542 (N1991,N1935,N1881);
nor U543 (N1995,N1938,N1886);
nor U544 (N1999,N1894,N1941);
nor U545 (N2000,N1941,N1891);
nor U546 (N2001,N1945,N1946);
nor U547 (N2004,N1902,N1947);
nor U548 (N2005,N1947,N1826);
nor U549 (N2006,N1905,N1951);
nor U550 (N2007,N1951,N1831);
nor U551 (N2008,N1908,N1955);
nor U552 (N2009,N1955,N1836);
nor U553 (N2010,N1911,N1959);
nor U554 (N2011,N1959,N1841);
nor U555 (N2012,N1914,N1963);
nor U556 (N2013,N1963,N1846);
nor U557 (N2014,N1917,N1967);
nor U558 (N2015,N1967,N1851);
nor U559 (N2016,N1920,N1971);
nor U560 (N2017,N1971,N1856);
nor U561 (N2018,N1923,N1975);
nor U562 (N2019,N1975,N1861);
nor U563 (N2020,N1926,N1979);
nor U564 (N2021,N1979,N1866);
nor U565 (N2022,N1929,N1983);
nor U566 (N2023,N1983,N1871);
nor U567 (N2024,N1932,N1987);
nor U568 (N2025,N1987,N1876);
nor U569 (N2026,N1935,N1991);
nor U570 (N2027,N1991,N1881);
nor U571 (N2028,N1938,N1995);
nor U572 (N2029,N1995,N1886);
nor U573 (N2030,N1999,N2000);
nor U574 (N2033,N2001,N1224);
nor U575 (N2037,N2004,N2005);
nor U576 (N2040,N2006,N2007);
nor U577 (N2043,N2008,N2009);
nor U578 (N2046,N2010,N2011);
nor U579 (N2049,N2012,N2013);
nor U580 (N2052,N2014,N2015);
nor U581 (N2055,N2016,N2017);
nor U582 (N2058,N2018,N2019);
nor U583 (N2061,N2020,N2021);
nor U584 (N2064,N2022,N2023);
nor U585 (N2067,N2024,N2025);
nor U586 (N2070,N2026,N2027);
nor U587 (N2073,N2028,N2029);
nor U588 (N2076,N2030,N1176);
nor U589 (N2080,N2001,N2033);
nor U590 (N2081,N2033,N1224);
nor U591 (N2082,N1897,N2033);
nor U592 (N2085,N2037,N552);
nor U593 (N2089,N2040,N600);
nor U594 (N2093,N2043,N648);
nor U595 (N2097,N2046,N696);
nor U596 (N2101,N2049,N744);
nor U597 (N2105,N2052,N792);
nor U598 (N2109,N2055,N840);
nor U599 (N2113,N2058,N888);
nor U600 (N2117,N2061,N936);
nor U601 (N2121,N2064,N984);
nor U602 (N2125,N2067,N1032);
nor U603 (N2129,N2070,N1080);
nor U604 (N2133,N2073,N1128);
nor U605 (N2137,N2030,N2076);
nor U606 (N2138,N2076,N1176);
nor U607 (N2139,N1941,N2076);
nor U608 (N2142,N2080,N2081);
nor U609 (N2145,N1272,N2082);
nor U610 (N2149,N2037,N2085);
nor U611 (N2150,N2085,N552);
nor U612 (N2151,N1947,N2085);
nor U613 (N2154,N2040,N2089);
nor U614 (N2155,N2089,N600);
nor U615 (N2156,N1951,N2089);
nor U616 (N2159,N2043,N2093);
nor U617 (N2160,N2093,N648);
nor U618 (N2161,N1955,N2093);
nor U619 (N2164,N2046,N2097);
nor U620 (N2165,N2097,N696);
nor U621 (N2166,N1959,N2097);
nor U622 (N2169,N2049,N2101);
nor U623 (N2170,N2101,N744);
nor U624 (N2171,N1963,N2101);
nor U625 (N2174,N2052,N2105);
nor U626 (N2175,N2105,N792);
nor U627 (N2176,N1967,N2105);
nor U628 (N2179,N2055,N2109);
nor U629 (N2180,N2109,N840);
nor U630 (N2181,N1971,N2109);
nor U631 (N2184,N2058,N2113);
nor U632 (N2185,N2113,N888);
nor U633 (N2186,N1975,N2113);
nor U634 (N2189,N2061,N2117);
nor U635 (N2190,N2117,N936);
nor U636 (N2191,N1979,N2117);
nor U637 (N2194,N2064,N2121);
nor U638 (N2195,N2121,N984);
nor U639 (N2196,N1983,N2121);
nor U640 (N2199,N2067,N2125);
nor U641 (N2200,N2125,N1032);
nor U642 (N2201,N1987,N2125);
nor U643 (N2204,N2070,N2129);
nor U644 (N2205,N2129,N1080);
nor U645 (N2206,N1991,N2129);
nor U646 (N2209,N2073,N2133);
nor U647 (N2210,N2133,N1128);
nor U648 (N2211,N1995,N2133);
nor U649 (N2214,N2137,N2138);
nor U650 (N2217,N2142,N2139);
nor U651 (N2221,N1272,N2145);
nor U652 (N2222,N2145,N2082);
nor U653 (N2223,N2149,N2150);
nor U654 (N2224,N2154,N2155);
nor U655 (N2227,N2159,N2160);
nor U656 (N2230,N2164,N2165);
nor U657 (N2233,N2169,N2170);
nor U658 (N2236,N2174,N2175);
nor U659 (N2239,N2179,N2180);
nor U660 (N2242,N2184,N2185);
nor U661 (N2245,N2189,N2190);
nor U662 (N2248,N2194,N2195);
nor U663 (N2251,N2199,N2200);
nor U664 (N2254,N2204,N2205);
nor U665 (N2257,N2209,N2210);
nor U666 (N2260,N2214,N2211);
nor U667 (N2264,N2142,N2217);
nor U668 (N2265,N2217,N2139);
nor U669 (N2266,N2221,N2222);
nor U670 (N2269,N2224,N2151);
nor U671 (N2273,N2227,N2156);
nor U672 (N2277,N2230,N2161);
nor U673 (N2281,N2233,N2166);
nor U674 (N2285,N2236,N2171);
nor U675 (N2289,N2239,N2176);
nor U676 (N2293,N2242,N2181);
nor U677 (N2297,N2245,N2186);
nor U678 (N2301,N2248,N2191);
nor U679 (N2305,N2251,N2196);
nor U680 (N2309,N2254,N2201);
nor U681 (N2313,N2257,N2206);
nor U682 (N2317,N2214,N2260);
nor U683 (N2318,N2260,N2211);
nor U684 (N2319,N2264,N2265);
nor U685 (N2322,N2266,N1227);
nor U686 (N2326,N2224,N2269);
nor U687 (N2327,N2269,N2151);
nor U688 (N2328,N2227,N2273);
nor U689 (N2329,N2273,N2156);
nor U690 (N2330,N2230,N2277);
nor U691 (N2331,N2277,N2161);
nor U692 (N2332,N2233,N2281);
nor U693 (N2333,N2281,N2166);
nor U694 (N2334,N2236,N2285);
nor U695 (N2335,N2285,N2171);
nor U696 (N2336,N2239,N2289);
nor U697 (N2337,N2289,N2176);
nor U698 (N2338,N2242,N2293);
nor U699 (N2339,N2293,N2181);
nor U700 (N2340,N2245,N2297);
nor U701 (N2341,N2297,N2186);
nor U702 (N2342,N2248,N2301);
nor U703 (N2343,N2301,N2191);
nor U704 (N2344,N2251,N2305);
nor U705 (N2345,N2305,N2196);
nor U706 (N2346,N2254,N2309);
nor U707 (N2347,N2309,N2201);
nor U708 (N2348,N2257,N2313);
nor U709 (N2349,N2313,N2206);
nor U710 (N2350,N2317,N2318);
nor U711 (N2353,N2319,N1179);
nor U712 (N2357,N2266,N2322);
nor U713 (N2358,N2322,N1227);
nor U714 (N2359,N2145,N2322);
nor U715 (N2362,N2326,N2327);
nor U716 (N2365,N2328,N2329);
nor U717 (N2368,N2330,N2331);
nor U718 (N2371,N2332,N2333);
nor U719 (N2374,N2334,N2335);
nor U720 (N2377,N2336,N2337);
nor U721 (N2380,N2338,N2339);
nor U722 (N2383,N2340,N2341);
nor U723 (N2386,N2342,N2343);
nor U724 (N2389,N2344,N2345);
nor U725 (N2392,N2346,N2347);
nor U726 (N2395,N2348,N2349);
nor U727 (N2398,N2350,N1131);
nor U728 (N2402,N2319,N2353);
nor U729 (N2403,N2353,N1179);
nor U730 (N2404,N2217,N2353);
nor U731 (N2407,N2357,N2358);
nor U732 (N2410,N1275,N2359);
nor U733 (N2414,N2362,N555);
nor U734 (N2418,N2365,N603);
nor U735 (N2422,N2368,N651);
nor U736 (N2426,N2371,N699);
nor U737 (N2430,N2374,N747);
nor U738 (N2434,N2377,N795);
nor U739 (N2438,N2380,N843);
nor U740 (N2442,N2383,N891);
nor U741 (N2446,N2386,N939);
nor U742 (N2450,N2389,N987);
nor U743 (N2454,N2392,N1035);
nor U744 (N2458,N2395,N1083);
nor U745 (N2462,N2350,N2398);
nor U746 (N2463,N2398,N1131);
nor U747 (N2464,N2260,N2398);
nor U748 (N2467,N2402,N2403);
nor U749 (N2470,N2407,N2404);
nor U750 (N2474,N1275,N2410);
nor U751 (N2475,N2410,N2359);
nor U752 (N2476,N2362,N2414);
nor U753 (N2477,N2414,N555);
nor U754 (N2478,N2269,N2414);
nor U755 (N2481,N2365,N2418);
nor U756 (N2482,N2418,N603);
nor U757 (N2483,N2273,N2418);
nor U758 (N2486,N2368,N2422);
nor U759 (N2487,N2422,N651);
nor U760 (N2488,N2277,N2422);
nor U761 (N2491,N2371,N2426);
nor U762 (N2492,N2426,N699);
nor U763 (N2493,N2281,N2426);
nor U764 (N2496,N2374,N2430);
nor U765 (N2497,N2430,N747);
nor U766 (N2498,N2285,N2430);
nor U767 (N2501,N2377,N2434);
nor U768 (N2502,N2434,N795);
nor U769 (N2503,N2289,N2434);
nor U770 (N2506,N2380,N2438);
nor U771 (N2507,N2438,N843);
nor U772 (N2508,N2293,N2438);
nor U773 (N2511,N2383,N2442);
nor U774 (N2512,N2442,N891);
nor U775 (N2513,N2297,N2442);
nor U776 (N2516,N2386,N2446);
nor U777 (N2517,N2446,N939);
nor U778 (N2518,N2301,N2446);
nor U779 (N2521,N2389,N2450);
nor U780 (N2522,N2450,N987);
nor U781 (N2523,N2305,N2450);
nor U782 (N2526,N2392,N2454);
nor U783 (N2527,N2454,N1035);
nor U784 (N2528,N2309,N2454);
nor U785 (N2531,N2395,N2458);
nor U786 (N2532,N2458,N1083);
nor U787 (N2533,N2313,N2458);
nor U788 (N2536,N2462,N2463);
nor U789 (N2539,N2467,N2464);
nor U790 (N2543,N2407,N2470);
nor U791 (N2544,N2470,N2404);
nor U792 (N2545,N2474,N2475);
nor U793 (N2548,N2476,N2477);
nor U794 (N2549,N2481,N2482);
nor U795 (N2552,N2486,N2487);
nor U796 (N2555,N2491,N2492);
nor U797 (N2558,N2496,N2497);
nor U798 (N2561,N2501,N2502);
nor U799 (N2564,N2506,N2507);
nor U800 (N2567,N2511,N2512);
nor U801 (N2570,N2516,N2517);
nor U802 (N2573,N2521,N2522);
nor U803 (N2576,N2526,N2527);
nor U804 (N2579,N2531,N2532);
nor U805 (N2582,N2536,N2533);
nor U806 (N2586,N2467,N2539);
nor U807 (N2587,N2539,N2464);
nor U808 (N2588,N2543,N2544);
nor U809 (N2591,N2545,N1230);
nor U810 (N2595,N2549,N2478);
nor U811 (N2599,N2552,N2483);
nor U812 (N2603,N2555,N2488);
nor U813 (N2607,N2558,N2493);
nor U814 (N2611,N2561,N2498);
nor U815 (N2615,N2564,N2503);
nor U816 (N2619,N2567,N2508);
nor U817 (N2623,N2570,N2513);
nor U818 (N2627,N2573,N2518);
nor U819 (N2631,N2576,N2523);
nor U820 (N2635,N2579,N2528);
nor U821 (N2639,N2536,N2582);
nor U822 (N2640,N2582,N2533);
nor U823 (N2641,N2586,N2587);
nor U824 (N2644,N2588,N1182);
nor U825 (N2648,N2545,N2591);
nor U826 (N2649,N2591,N1230);
nor U827 (N2650,N2410,N2591);
nor U828 (N2653,N2549,N2595);
nor U829 (N2654,N2595,N2478);
nor U830 (N2655,N2552,N2599);
nor U831 (N2656,N2599,N2483);
nor U832 (N2657,N2555,N2603);
nor U833 (N2658,N2603,N2488);
nor U834 (N2659,N2558,N2607);
nor U835 (N2660,N2607,N2493);
nor U836 (N2661,N2561,N2611);
nor U837 (N2662,N2611,N2498);
nor U838 (N2663,N2564,N2615);
nor U839 (N2664,N2615,N2503);
nor U840 (N2665,N2567,N2619);
nor U841 (N2666,N2619,N2508);
nor U842 (N2667,N2570,N2623);
nor U843 (N2668,N2623,N2513);
nor U844 (N2669,N2573,N2627);
nor U845 (N2670,N2627,N2518);
nor U846 (N2671,N2576,N2631);
nor U847 (N2672,N2631,N2523);
nor U848 (N2673,N2579,N2635);
nor U849 (N2674,N2635,N2528);
nor U850 (N2675,N2639,N2640);
nor U851 (N2678,N2641,N1134);
nor U852 (N2682,N2588,N2644);
nor U853 (N2683,N2644,N1182);
nor U854 (N2684,N2470,N2644);
nor U855 (N2687,N2648,N2649);
nor U856 (N2690,N1278,N2650);
nor U857 (N2694,N2653,N2654);
nor U858 (N2697,N2655,N2656);
nor U859 (N2700,N2657,N2658);
nor U860 (N2703,N2659,N2660);
nor U861 (N2706,N2661,N2662);
nor U862 (N2709,N2663,N2664);
nor U863 (N2712,N2665,N2666);
nor U864 (N2715,N2667,N2668);
nor U865 (N2718,N2669,N2670);
nor U866 (N2721,N2671,N2672);
nor U867 (N2724,N2673,N2674);
nor U868 (N2727,N2675,N1086);
nor U869 (N2731,N2641,N2678);
nor U870 (N2732,N2678,N1134);
nor U871 (N2733,N2539,N2678);
nor U872 (N2736,N2682,N2683);
nor U873 (N2739,N2687,N2684);
nor U874 (N2743,N1278,N2690);
nor U875 (N2744,N2690,N2650);
nor U876 (N2745,N2694,N558);
nor U877 (N2749,N2697,N606);
nor U878 (N2753,N2700,N654);
nor U879 (N2757,N2703,N702);
nor U880 (N2761,N2706,N750);
nor U881 (N2765,N2709,N798);
nor U882 (N2769,N2712,N846);
nor U883 (N2773,N2715,N894);
nor U884 (N2777,N2718,N942);
nor U885 (N2781,N2721,N990);
nor U886 (N2785,N2724,N1038);
nor U887 (N2789,N2675,N2727);
nor U888 (N2790,N2727,N1086);
nor U889 (N2791,N2582,N2727);
nor U890 (N2794,N2731,N2732);
nor U891 (N2797,N2736,N2733);
nor U892 (N2801,N2687,N2739);
nor U893 (N2802,N2739,N2684);
nor U894 (N2803,N2743,N2744);
nor U895 (N2806,N2694,N2745);
nor U896 (N2807,N2745,N558);
nor U897 (N2808,N2595,N2745);
nor U898 (N2811,N2697,N2749);
nor U899 (N2812,N2749,N606);
nor U900 (N2813,N2599,N2749);
nor U901 (N2816,N2700,N2753);
nor U902 (N2817,N2753,N654);
nor U903 (N2818,N2603,N2753);
nor U904 (N2821,N2703,N2757);
nor U905 (N2822,N2757,N702);
nor U906 (N2823,N2607,N2757);
nor U907 (N2826,N2706,N2761);
nor U908 (N2827,N2761,N750);
nor U909 (N2828,N2611,N2761);
nor U910 (N2831,N2709,N2765);
nor U911 (N2832,N2765,N798);
nor U912 (N2833,N2615,N2765);
nor U913 (N2836,N2712,N2769);
nor U914 (N2837,N2769,N846);
nor U915 (N2838,N2619,N2769);
nor U916 (N2841,N2715,N2773);
nor U917 (N2842,N2773,N894);
nor U918 (N2843,N2623,N2773);
nor U919 (N2846,N2718,N2777);
nor U920 (N2847,N2777,N942);
nor U921 (N2848,N2627,N2777);
nor U922 (N2851,N2721,N2781);
nor U923 (N2852,N2781,N990);
nor U924 (N2853,N2631,N2781);
nor U925 (N2856,N2724,N2785);
nor U926 (N2857,N2785,N1038);
nor U927 (N2858,N2635,N2785);
nor U928 (N2861,N2789,N2790);
nor U929 (N2864,N2794,N2791);
nor U930 (N2868,N2736,N2797);
nor U931 (N2869,N2797,N2733);
nor U932 (N2870,N2801,N2802);
nor U933 (N2873,N2803,N1233);
nor U934 (N2877,N2806,N2807);
nor U935 (N2878,N2811,N2812);
nor U936 (N2881,N2816,N2817);
nor U937 (N2884,N2821,N2822);
nor U938 (N2887,N2826,N2827);
nor U939 (N2890,N2831,N2832);
nor U940 (N2893,N2836,N2837);
nor U941 (N2896,N2841,N2842);
nor U942 (N2899,N2846,N2847);
nor U943 (N2902,N2851,N2852);
nor U944 (N2905,N2856,N2857);
nor U945 (N2908,N2861,N2858);
nor U946 (N2912,N2794,N2864);
nor U947 (N2913,N2864,N2791);
nor U948 (N2914,N2868,N2869);
nor U949 (N2917,N2870,N1185);
nor U950 (N2921,N2803,N2873);
nor U951 (N2922,N2873,N1233);
nor U952 (N2923,N2690,N2873);
nor U953 (N2926,N2878,N2808);
nor U954 (N2930,N2881,N2813);
nor U955 (N2934,N2884,N2818);
nor U956 (N2938,N2887,N2823);
nor U957 (N2942,N2890,N2828);
nor U958 (N2946,N2893,N2833);
nor U959 (N2950,N2896,N2838);
nor U960 (N2954,N2899,N2843);
nor U961 (N2958,N2902,N2848);
nor U962 (N2962,N2905,N2853);
nor U963 (N2966,N2861,N2908);
nor U964 (N2967,N2908,N2858);
nor U965 (N2968,N2912,N2913);
nor U966 (N2971,N2914,N1137);
nor U967 (N2975,N2870,N2917);
nor U968 (N2976,N2917,N1185);
nor U969 (N2977,N2739,N2917);
nor U970 (N2980,N2921,N2922);
nor U971 (N2983,N1281,N2923);
nor U972 (N2987,N2878,N2926);
nor U973 (N2988,N2926,N2808);
nor U974 (N2989,N2881,N2930);
nor U975 (N2990,N2930,N2813);
nor U976 (N2991,N2884,N2934);
nor U977 (N2992,N2934,N2818);
nor U978 (N2993,N2887,N2938);
nor U979 (N2994,N2938,N2823);
nor U980 (N2995,N2890,N2942);
nor U981 (N2996,N2942,N2828);
nor U982 (N2997,N2893,N2946);
nor U983 (N2998,N2946,N2833);
nor U984 (N2999,N2896,N2950);
nor U985 (N3000,N2950,N2838);
nor U986 (N3001,N2899,N2954);
nor U987 (N3002,N2954,N2843);
nor U988 (N3003,N2902,N2958);
nor U989 (N3004,N2958,N2848);
nor U990 (N3005,N2905,N2962);
nor U991 (N3006,N2962,N2853);
nor U992 (N3007,N2966,N2967);
nor U993 (N3010,N2968,N1089);
nor U994 (N3014,N2914,N2971);
nor U995 (N3015,N2971,N1137);
nor U996 (N3016,N2797,N2971);
nor U997 (N3019,N2975,N2976);
nor U998 (N3022,N2980,N2977);
nor U999 (N3026,N1281,N2983);
nor U1000 (N3027,N2983,N2923);
nor U1001 (N3028,N2987,N2988);
nor U1002 (N3031,N2989,N2990);
nor U1003 (N3034,N2991,N2992);
nor U1004 (N3037,N2993,N2994);
nor U1005 (N3040,N2995,N2996);
nor U1006 (N3043,N2997,N2998);
nor U1007 (N3046,N2999,N3000);
nor U1008 (N3049,N3001,N3002);
nor U1009 (N3052,N3003,N3004);
nor U1010 (N3055,N3005,N3006);
nor U1011 (N3058,N3007,N1041);
nor U1012 (N3062,N2968,N3010);
nor U1013 (N3063,N3010,N1089);
nor U1014 (N3064,N2864,N3010);
nor U1015 (N3067,N3014,N3015);
nor U1016 (N3070,N3019,N3016);
nor U1017 (N3074,N2980,N3022);
nor U1018 (N3075,N3022,N2977);
nor U1019 (N3076,N3026,N3027);
nor U1020 (N3079,N3028,N561);
nor U1021 (N3083,N3031,N609);
nor U1022 (N3087,N3034,N657);
nor U1023 (N3091,N3037,N705);
nor U1024 (N3095,N3040,N753);
nor U1025 (N3099,N3043,N801);
nor U1026 (N3103,N3046,N849);
nor U1027 (N3107,N3049,N897);
nor U1028 (N3111,N3052,N945);
nor U1029 (N3115,N3055,N993);
nor U1030 (N3119,N3007,N3058);
nor U1031 (N3120,N3058,N1041);
nor U1032 (N3121,N2908,N3058);
nor U1033 (N3124,N3062,N3063);
nor U1034 (N3127,N3067,N3064);
nor U1035 (N3131,N3019,N3070);
nor U1036 (N3132,N3070,N3016);
nor U1037 (N3133,N3074,N3075);
nor U1038 (N3136,N3076,N1236);
nor U1039 (N3140,N3028,N3079);
nor U1040 (N3141,N3079,N561);
nor U1041 (N3142,N2926,N3079);
nor U1042 (N3145,N3031,N3083);
nor U1043 (N3146,N3083,N609);
nor U1044 (N3147,N2930,N3083);
nor U1045 (N3150,N3034,N3087);
nor U1046 (N3151,N3087,N657);
nor U1047 (N3152,N2934,N3087);
nor U1048 (N3155,N3037,N3091);
nor U1049 (N3156,N3091,N705);
nor U1050 (N3157,N2938,N3091);
nor U1051 (N3160,N3040,N3095);
nor U1052 (N3161,N3095,N753);
nor U1053 (N3162,N2942,N3095);
nor U1054 (N3165,N3043,N3099);
nor U1055 (N3166,N3099,N801);
nor U1056 (N3167,N2946,N3099);
nor U1057 (N3170,N3046,N3103);
nor U1058 (N3171,N3103,N849);
nor U1059 (N3172,N2950,N3103);
nor U1060 (N3175,N3049,N3107);
nor U1061 (N3176,N3107,N897);
nor U1062 (N3177,N2954,N3107);
nor U1063 (N3180,N3052,N3111);
nor U1064 (N3181,N3111,N945);
nor U1065 (N3182,N2958,N3111);
nor U1066 (N3185,N3055,N3115);
nor U1067 (N3186,N3115,N993);
nor U1068 (N3187,N2962,N3115);
nor U1069 (N3190,N3119,N3120);
nor U1070 (N3193,N3124,N3121);
nor U1071 (N3197,N3067,N3127);
nor U1072 (N3198,N3127,N3064);
nor U1073 (N3199,N3131,N3132);
nor U1074 (N3202,N3133,N1188);
nor U1075 (N3206,N3076,N3136);
nor U1076 (N3207,N3136,N1236);
nor U1077 (N3208,N2983,N3136);
nor U1078 (N3211,N3140,N3141);
nor U1079 (N3212,N3145,N3146);
nor U1080 (N3215,N3150,N3151);
nor U1081 (N3218,N3155,N3156);
nor U1082 (N3221,N3160,N3161);
nor U1083 (N3224,N3165,N3166);
nor U1084 (N3227,N3170,N3171);
nor U1085 (N3230,N3175,N3176);
nor U1086 (N3233,N3180,N3181);
nor U1087 (N3236,N3185,N3186);
nor U1088 (N3239,N3190,N3187);
nor U1089 (N3243,N3124,N3193);
nor U1090 (N3244,N3193,N3121);
nor U1091 (N3245,N3197,N3198);
nor U1092 (N3248,N3199,N1140);
nor U1093 (N3252,N3133,N3202);
nor U1094 (N3253,N3202,N1188);
nor U1095 (N3254,N3022,N3202);
nor U1096 (N3257,N3206,N3207);
nor U1097 (N3260,N1284,N3208);
nor U1098 (N3264,N3212,N3142);
nor U1099 (N3268,N3215,N3147);
nor U1100 (N3272,N3218,N3152);
nor U1101 (N3276,N3221,N3157);
nor U1102 (N3280,N3224,N3162);
nor U1103 (N3284,N3227,N3167);
nor U1104 (N3288,N3230,N3172);
nor U1105 (N3292,N3233,N3177);
nor U1106 (N3296,N3236,N3182);
nor U1107 (N3300,N3190,N3239);
nor U1108 (N3301,N3239,N3187);
nor U1109 (N3302,N3243,N3244);
nor U1110 (N3305,N3245,N1092);
nor U1111 (N3309,N3199,N3248);
nor U1112 (N3310,N3248,N1140);
nor U1113 (N3311,N3070,N3248);
nor U1114 (N3314,N3252,N3253);
nor U1115 (N3317,N3257,N3254);
nor U1116 (N3321,N1284,N3260);
nor U1117 (N3322,N3260,N3208);
nor U1118 (N3323,N3212,N3264);
nor U1119 (N3324,N3264,N3142);
nor U1120 (N3325,N3215,N3268);
nor U1121 (N3326,N3268,N3147);
nor U1122 (N3327,N3218,N3272);
nor U1123 (N3328,N3272,N3152);
nor U1124 (N3329,N3221,N3276);
nor U1125 (N3330,N3276,N3157);
nor U1126 (N3331,N3224,N3280);
nor U1127 (N3332,N3280,N3162);
nor U1128 (N3333,N3227,N3284);
nor U1129 (N3334,N3284,N3167);
nor U1130 (N3335,N3230,N3288);
nor U1131 (N3336,N3288,N3172);
nor U1132 (N3337,N3233,N3292);
nor U1133 (N3338,N3292,N3177);
nor U1134 (N3339,N3236,N3296);
nor U1135 (N3340,N3296,N3182);
nor U1136 (N3341,N3300,N3301);
nor U1137 (N3344,N3302,N1044);
nor U1138 (N3348,N3245,N3305);
nor U1139 (N3349,N3305,N1092);
nor U1140 (N3350,N3127,N3305);
nor U1141 (N3353,N3309,N3310);
nor U1142 (N3356,N3314,N3311);
nor U1143 (N3360,N3257,N3317);
nor U1144 (N3361,N3317,N3254);
nor U1145 (N3362,N3321,N3322);
nor U1146 (N3365,N3323,N3324);
nor U1147 (N3368,N3325,N3326);
nor U1148 (N3371,N3327,N3328);
nor U1149 (N3374,N3329,N3330);
nor U1150 (N3377,N3331,N3332);
nor U1151 (N3380,N3333,N3334);
nor U1152 (N3383,N3335,N3336);
nor U1153 (N3386,N3337,N3338);
nor U1154 (N3389,N3339,N3340);
nor U1155 (N3392,N3341,N996);
nor U1156 (N3396,N3302,N3344);
nor U1157 (N3397,N3344,N1044);
nor U1158 (N3398,N3193,N3344);
nor U1159 (N3401,N3348,N3349);
nor U1160 (N3404,N3353,N3350);
nor U1161 (N3408,N3314,N3356);
nor U1162 (N3409,N3356,N3311);
nor U1163 (N3410,N3360,N3361);
nor U1164 (N3413,N3362,N1239);
nor U1165 (N3417,N3365,N564);
nor U1166 (N3421,N3368,N612);
nor U1167 (N3425,N3371,N660);
nor U1168 (N3429,N3374,N708);
nor U1169 (N3433,N3377,N756);
nor U1170 (N3437,N3380,N804);
nor U1171 (N3441,N3383,N852);
nor U1172 (N3445,N3386,N900);
nor U1173 (N3449,N3389,N948);
nor U1174 (N3453,N3341,N3392);
nor U1175 (N3454,N3392,N996);
nor U1176 (N3455,N3239,N3392);
nor U1177 (N3458,N3396,N3397);
nor U1178 (N3461,N3401,N3398);
nor U1179 (N3465,N3353,N3404);
nor U1180 (N3466,N3404,N3350);
nor U1181 (N3467,N3408,N3409);
nor U1182 (N3470,N3410,N1191);
nor U1183 (N3474,N3362,N3413);
nor U1184 (N3475,N3413,N1239);
nor U1185 (N3476,N3260,N3413);
nor U1186 (N3479,N3365,N3417);
nor U1187 (N3480,N3417,N564);
nor U1188 (N3481,N3264,N3417);
nor U1189 (N3484,N3368,N3421);
nor U1190 (N3485,N3421,N612);
nor U1191 (N3486,N3268,N3421);
nor U1192 (N3489,N3371,N3425);
nor U1193 (N3490,N3425,N660);
nor U1194 (N3491,N3272,N3425);
nor U1195 (N3494,N3374,N3429);
nor U1196 (N3495,N3429,N708);
nor U1197 (N3496,N3276,N3429);
nor U1198 (N3499,N3377,N3433);
nor U1199 (N3500,N3433,N756);
nor U1200 (N3501,N3280,N3433);
nor U1201 (N3504,N3380,N3437);
nor U1202 (N3505,N3437,N804);
nor U1203 (N3506,N3284,N3437);
nor U1204 (N3509,N3383,N3441);
nor U1205 (N3510,N3441,N852);
nor U1206 (N3511,N3288,N3441);
nor U1207 (N3514,N3386,N3445);
nor U1208 (N3515,N3445,N900);
nor U1209 (N3516,N3292,N3445);
nor U1210 (N3519,N3389,N3449);
nor U1211 (N3520,N3449,N948);
nor U1212 (N3521,N3296,N3449);
nor U1213 (N3524,N3453,N3454);
nor U1214 (N3527,N3458,N3455);
nor U1215 (N3531,N3401,N3461);
nor U1216 (N3532,N3461,N3398);
nor U1217 (N3533,N3465,N3466);
nor U1218 (N3536,N3467,N1143);
nor U1219 (N3540,N3410,N3470);
nor U1220 (N3541,N3470,N1191);
nor U1221 (N3542,N3317,N3470);
nor U1222 (N3545,N3474,N3475);
nor U1223 (N3548,N1287,N3476);
nor U1224 (N3552,N3479,N3480);
nor U1225 (N3553,N3484,N3485);
nor U1226 (N3556,N3489,N3490);
nor U1227 (N3559,N3494,N3495);
nor U1228 (N3562,N3499,N3500);
nor U1229 (N3565,N3504,N3505);
nor U1230 (N3568,N3509,N3510);
nor U1231 (N3571,N3514,N3515);
nor U1232 (N3574,N3519,N3520);
nor U1233 (N3577,N3524,N3521);
nor U1234 (N3581,N3458,N3527);
nor U1235 (N3582,N3527,N3455);
nor U1236 (N3583,N3531,N3532);
nor U1237 (N3586,N3533,N1095);
nor U1238 (N3590,N3467,N3536);
nor U1239 (N3591,N3536,N1143);
nor U1240 (N3592,N3356,N3536);
nor U1241 (N3595,N3540,N3541);
nor U1242 (N3598,N3545,N3542);
nor U1243 (N3602,N1287,N3548);
nor U1244 (N3603,N3548,N3476);
nor U1245 (N3604,N3553,N3481);
nor U1246 (N3608,N3556,N3486);
nor U1247 (N3612,N3559,N3491);
nor U1248 (N3616,N3562,N3496);
nor U1249 (N3620,N3565,N3501);
nor U1250 (N3624,N3568,N3506);
nor U1251 (N3628,N3571,N3511);
nor U1252 (N3632,N3574,N3516);
nor U1253 (N3636,N3524,N3577);
nor U1254 (N3637,N3577,N3521);
nor U1255 (N3638,N3581,N3582);
nor U1256 (N3641,N3583,N1047);
nor U1257 (N3645,N3533,N3586);
nor U1258 (N3646,N3586,N1095);
nor U1259 (N3647,N3404,N3586);
nor U1260 (N3650,N3590,N3591);
nor U1261 (N3653,N3595,N3592);
nor U1262 (N3657,N3545,N3598);
nor U1263 (N3658,N3598,N3542);
nor U1264 (N3659,N3602,N3603);
nor U1265 (N3662,N3553,N3604);
nor U1266 (N3663,N3604,N3481);
nor U1267 (N3664,N3556,N3608);
nor U1268 (N3665,N3608,N3486);
nor U1269 (N3666,N3559,N3612);
nor U1270 (N3667,N3612,N3491);
nor U1271 (N3668,N3562,N3616);
nor U1272 (N3669,N3616,N3496);
nor U1273 (N3670,N3565,N3620);
nor U1274 (N3671,N3620,N3501);
nor U1275 (N3672,N3568,N3624);
nor U1276 (N3673,N3624,N3506);
nor U1277 (N3674,N3571,N3628);
nor U1278 (N3675,N3628,N3511);
nor U1279 (N3676,N3574,N3632);
nor U1280 (N3677,N3632,N3516);
nor U1281 (N3678,N3636,N3637);
nor U1282 (N3681,N3638,N999);
nor U1283 (N3685,N3583,N3641);
nor U1284 (N3686,N3641,N1047);
nor U1285 (N3687,N3461,N3641);
nor U1286 (N3690,N3645,N3646);
nor U1287 (N3693,N3650,N3647);
nor U1288 (N3697,N3595,N3653);
nor U1289 (N3698,N3653,N3592);
nor U1290 (N3699,N3657,N3658);
nor U1291 (N3702,N3659,N1242);
nor U1292 (N3706,N3662,N3663);
nor U1293 (N3709,N3664,N3665);
nor U1294 (N3712,N3666,N3667);
nor U1295 (N3715,N3668,N3669);
nor U1296 (N3718,N3670,N3671);
nor U1297 (N3721,N3672,N3673);
nor U1298 (N3724,N3674,N3675);
nor U1299 (N3727,N3676,N3677);
nor U1300 (N3730,N3678,N951);
nor U1301 (N3734,N3638,N3681);
nor U1302 (N3735,N3681,N999);
nor U1303 (N3736,N3527,N3681);
nor U1304 (N3739,N3685,N3686);
nor U1305 (N3742,N3690,N3687);
nor U1306 (N3746,N3650,N3693);
nor U1307 (N3747,N3693,N3647);
nor U1308 (N3748,N3697,N3698);
nor U1309 (N3751,N3699,N1194);
nor U1310 (N3755,N3659,N3702);
nor U1311 (N3756,N3702,N1242);
nor U1312 (N3757,N3548,N3702);
nor U1313 (N3760,N3706,N567);
nor U1314 (N3764,N3709,N615);
nor U1315 (N3768,N3712,N663);
nor U1316 (N3772,N3715,N711);
nor U1317 (N3776,N3718,N759);
nor U1318 (N3780,N3721,N807);
nor U1319 (N3784,N3724,N855);
nor U1320 (N3788,N3727,N903);
nor U1321 (N3792,N3678,N3730);
nor U1322 (N3793,N3730,N951);
nor U1323 (N3794,N3577,N3730);
nor U1324 (N3797,N3734,N3735);
nor U1325 (N3800,N3739,N3736);
nor U1326 (N3804,N3690,N3742);
nor U1327 (N3805,N3742,N3687);
nor U1328 (N3806,N3746,N3747);
nor U1329 (N3809,N3748,N1146);
nor U1330 (N3813,N3699,N3751);
nor U1331 (N3814,N3751,N1194);
nor U1332 (N3815,N3598,N3751);
nor U1333 (N3818,N3755,N3756);
nor U1334 (N3821,N1290,N3757);
nor U1335 (N3825,N3706,N3760);
nor U1336 (N3826,N3760,N567);
nor U1337 (N3827,N3604,N3760);
nor U1338 (N3830,N3709,N3764);
nor U1339 (N3831,N3764,N615);
nor U1340 (N3832,N3608,N3764);
nor U1341 (N3835,N3712,N3768);
nor U1342 (N3836,N3768,N663);
nor U1343 (N3837,N3612,N3768);
nor U1344 (N3840,N3715,N3772);
nor U1345 (N3841,N3772,N711);
nor U1346 (N3842,N3616,N3772);
nor U1347 (N3845,N3718,N3776);
nor U1348 (N3846,N3776,N759);
nor U1349 (N3847,N3620,N3776);
nor U1350 (N3850,N3721,N3780);
nor U1351 (N3851,N3780,N807);
nor U1352 (N3852,N3624,N3780);
nor U1353 (N3855,N3724,N3784);
nor U1354 (N3856,N3784,N855);
nor U1355 (N3857,N3628,N3784);
nor U1356 (N3860,N3727,N3788);
nor U1357 (N3861,N3788,N903);
nor U1358 (N3862,N3632,N3788);
nor U1359 (N3865,N3792,N3793);
nor U1360 (N3868,N3797,N3794);
nor U1361 (N3872,N3739,N3800);
nor U1362 (N3873,N3800,N3736);
nor U1363 (N3874,N3804,N3805);
nor U1364 (N3877,N3806,N1098);
nor U1365 (N3881,N3748,N3809);
nor U1366 (N3882,N3809,N1146);
nor U1367 (N3883,N3653,N3809);
nor U1368 (N3886,N3813,N3814);
nor U1369 (N3889,N3818,N3815);
nor U1370 (N3893,N1290,N3821);
nor U1371 (N3894,N3821,N3757);
nor U1372 (N3895,N3825,N3826);
nor U1373 (N3896,N3830,N3831);
nor U1374 (N3899,N3835,N3836);
nor U1375 (N3902,N3840,N3841);
nor U1376 (N3905,N3845,N3846);
nor U1377 (N3908,N3850,N3851);
nor U1378 (N3911,N3855,N3856);
nor U1379 (N3914,N3860,N3861);
nor U1380 (N3917,N3865,N3862);
nor U1381 (N3921,N3797,N3868);
nor U1382 (N3922,N3868,N3794);
nor U1383 (N3923,N3872,N3873);
nor U1384 (N3926,N3874,N1050);
nor U1385 (N3930,N3806,N3877);
nor U1386 (N3931,N3877,N1098);
nor U1387 (N3932,N3693,N3877);
nor U1388 (N3935,N3881,N3882);
nor U1389 (N3938,N3886,N3883);
nor U1390 (N3942,N3818,N3889);
nor U1391 (N3943,N3889,N3815);
nor U1392 (N3944,N3893,N3894);
nor U1393 (N3947,N3896,N3827);
nor U1394 (N3951,N3899,N3832);
nor U1395 (N3955,N3902,N3837);
nor U1396 (N3959,N3905,N3842);
nor U1397 (N3963,N3908,N3847);
nor U1398 (N3967,N3911,N3852);
nor U1399 (N3971,N3914,N3857);
nor U1400 (N3975,N3865,N3917);
nor U1401 (N3976,N3917,N3862);
nor U1402 (N3977,N3921,N3922);
nor U1403 (N3980,N3923,N1002);
nor U1404 (N3984,N3874,N3926);
nor U1405 (N3985,N3926,N1050);
nor U1406 (N3986,N3742,N3926);
nor U1407 (N3989,N3930,N3931);
nor U1408 (N3992,N3935,N3932);
nor U1409 (N3996,N3886,N3938);
nor U1410 (N3997,N3938,N3883);
nor U1411 (N3998,N3942,N3943);
nor U1412 (N4001,N3944,N1245);
nor U1413 (N4005,N3896,N3947);
nor U1414 (N4006,N3947,N3827);
nor U1415 (N4007,N3899,N3951);
nor U1416 (N4008,N3951,N3832);
nor U1417 (N4009,N3902,N3955);
nor U1418 (N4010,N3955,N3837);
nor U1419 (N4011,N3905,N3959);
nor U1420 (N4012,N3959,N3842);
nor U1421 (N4013,N3908,N3963);
nor U1422 (N4014,N3963,N3847);
nor U1423 (N4015,N3911,N3967);
nor U1424 (N4016,N3967,N3852);
nor U1425 (N4017,N3914,N3971);
nor U1426 (N4018,N3971,N3857);
nor U1427 (N4019,N3975,N3976);
nor U1428 (N4022,N3977,N954);
nor U1429 (N4026,N3923,N3980);
nor U1430 (N4027,N3980,N1002);
nor U1431 (N4028,N3800,N3980);
nor U1432 (N4031,N3984,N3985);
nor U1433 (N4034,N3989,N3986);
nor U1434 (N4038,N3935,N3992);
nor U1435 (N4039,N3992,N3932);
nor U1436 (N4040,N3996,N3997);
nor U1437 (N4043,N3998,N1197);
nor U1438 (N4047,N3944,N4001);
nor U1439 (N4048,N4001,N1245);
nor U1440 (N4049,N3821,N4001);
nor U1441 (N4052,N4005,N4006);
nor U1442 (N4055,N4007,N4008);
nor U1443 (N4058,N4009,N4010);
nor U1444 (N4061,N4011,N4012);
nor U1445 (N4064,N4013,N4014);
nor U1446 (N4067,N4015,N4016);
nor U1447 (N4070,N4017,N4018);
nor U1448 (N4073,N4019,N906);
nor U1449 (N4077,N3977,N4022);
nor U1450 (N4078,N4022,N954);
nor U1451 (N4079,N3868,N4022);
nor U1452 (N4082,N4026,N4027);
nor U1453 (N4085,N4031,N4028);
nor U1454 (N4089,N3989,N4034);
nor U1455 (N4090,N4034,N3986);
nor U1456 (N4091,N4038,N4039);
nor U1457 (N4094,N4040,N1149);
nor U1458 (N4098,N3998,N4043);
nor U1459 (N4099,N4043,N1197);
nor U1460 (N4100,N3889,N4043);
nor U1461 (N4103,N4047,N4048);
nor U1462 (N4106,N1293,N4049);
nor U1463 (N4110,N4052,N570);
nor U1464 (N4114,N4055,N618);
nor U1465 (N4118,N4058,N666);
nor U1466 (N4122,N4061,N714);
nor U1467 (N4126,N4064,N762);
nor U1468 (N4130,N4067,N810);
nor U1469 (N4134,N4070,N858);
nor U1470 (N4138,N4019,N4073);
nor U1471 (N4139,N4073,N906);
nor U1472 (N4140,N3917,N4073);
nor U1473 (N4143,N4077,N4078);
nor U1474 (N4146,N4082,N4079);
nor U1475 (N4150,N4031,N4085);
nor U1476 (N4151,N4085,N4028);
nor U1477 (N4152,N4089,N4090);
nor U1478 (N4155,N4091,N1101);
nor U1479 (N4159,N4040,N4094);
nor U1480 (N4160,N4094,N1149);
nor U1481 (N4161,N3938,N4094);
nor U1482 (N4164,N4098,N4099);
nor U1483 (N4167,N4103,N4100);
nor U1484 (N4171,N1293,N4106);
nor U1485 (N4172,N4106,N4049);
nor U1486 (N4173,N4052,N4110);
nor U1487 (N4174,N4110,N570);
nor U1488 (N4175,N3947,N4110);
nor U1489 (N4178,N4055,N4114);
nor U1490 (N4179,N4114,N618);
nor U1491 (N4180,N3951,N4114);
nor U1492 (N4183,N4058,N4118);
nor U1493 (N4184,N4118,N666);
nor U1494 (N4185,N3955,N4118);
nor U1495 (N4188,N4061,N4122);
nor U1496 (N4189,N4122,N714);
nor U1497 (N4190,N3959,N4122);
nor U1498 (N4193,N4064,N4126);
nor U1499 (N4194,N4126,N762);
nor U1500 (N4195,N3963,N4126);
nor U1501 (N4198,N4067,N4130);
nor U1502 (N4199,N4130,N810);
nor U1503 (N4200,N3967,N4130);
nor U1504 (N4203,N4070,N4134);
nor U1505 (N4204,N4134,N858);
nor U1506 (N4205,N3971,N4134);
nor U1507 (N4208,N4138,N4139);
nor U1508 (N4211,N4143,N4140);
nor U1509 (N4215,N4082,N4146);
nor U1510 (N4216,N4146,N4079);
nor U1511 (N4217,N4150,N4151);
nor U1512 (N4220,N4152,N1053);
nor U1513 (N4224,N4091,N4155);
nor U1514 (N4225,N4155,N1101);
nor U1515 (N4226,N3992,N4155);
nor U1516 (N4229,N4159,N4160);
nor U1517 (N4232,N4164,N4161);
nor U1518 (N4236,N4103,N4167);
nor U1519 (N4237,N4167,N4100);
nor U1520 (N4238,N4171,N4172);
nor U1521 (N4241,N4173,N4174);
nor U1522 (N4242,N4178,N4179);
nor U1523 (N4245,N4183,N4184);
nor U1524 (N4248,N4188,N4189);
nor U1525 (N4251,N4193,N4194);
nor U1526 (N4254,N4198,N4199);
nor U1527 (N4257,N4203,N4204);
nor U1528 (N4260,N4208,N4205);
nor U1529 (N4264,N4143,N4211);
nor U1530 (N4265,N4211,N4140);
nor U1531 (N4266,N4215,N4216);
nor U1532 (N4269,N4217,N1005);
nor U1533 (N4273,N4152,N4220);
nor U1534 (N4274,N4220,N1053);
nor U1535 (N4275,N4034,N4220);
nor U1536 (N4278,N4224,N4225);
nor U1537 (N4281,N4229,N4226);
nor U1538 (N4285,N4164,N4232);
nor U1539 (N4286,N4232,N4161);
nor U1540 (N4287,N4236,N4237);
nor U1541 (N4290,N4238,N1248);
nor U1542 (N4294,N4242,N4175);
nor U1543 (N4298,N4245,N4180);
nor U1544 (N4302,N4248,N4185);
nor U1545 (N4306,N4251,N4190);
nor U1546 (N4310,N4254,N4195);
nor U1547 (N4314,N4257,N4200);
nor U1548 (N4318,N4208,N4260);
nor U1549 (N4319,N4260,N4205);
nor U1550 (N4320,N4264,N4265);
nor U1551 (N4323,N4266,N957);
nor U1552 (N4327,N4217,N4269);
nor U1553 (N4328,N4269,N1005);
nor U1554 (N4329,N4085,N4269);
nor U1555 (N4332,N4273,N4274);
nor U1556 (N4335,N4278,N4275);
nor U1557 (N4339,N4229,N4281);
nor U1558 (N4340,N4281,N4226);
nor U1559 (N4341,N4285,N4286);
nor U1560 (N4344,N4287,N1200);
nor U1561 (N4348,N4238,N4290);
nor U1562 (N4349,N4290,N1248);
nor U1563 (N4350,N4106,N4290);
nor U1564 (N4353,N4242,N4294);
nor U1565 (N4354,N4294,N4175);
nor U1566 (N4355,N4245,N4298);
nor U1567 (N4356,N4298,N4180);
nor U1568 (N4357,N4248,N4302);
nor U1569 (N4358,N4302,N4185);
nor U1570 (N4359,N4251,N4306);
nor U1571 (N4360,N4306,N4190);
nor U1572 (N4361,N4254,N4310);
nor U1573 (N4362,N4310,N4195);
nor U1574 (N4363,N4257,N4314);
nor U1575 (N4364,N4314,N4200);
nor U1576 (N4365,N4318,N4319);
nor U1577 (N4368,N4320,N909);
nor U1578 (N4372,N4266,N4323);
nor U1579 (N4373,N4323,N957);
nor U1580 (N4374,N4146,N4323);
nor U1581 (N4377,N4327,N4328);
nor U1582 (N4380,N4332,N4329);
nor U1583 (N4384,N4278,N4335);
nor U1584 (N4385,N4335,N4275);
nor U1585 (N4386,N4339,N4340);
nor U1586 (N4389,N4341,N1152);
nor U1587 (N4393,N4287,N4344);
nor U1588 (N4394,N4344,N1200);
nor U1589 (N4395,N4167,N4344);
nor U1590 (N4398,N4348,N4349);
nor U1591 (N4401,N1296,N4350);
nor U1592 (N4405,N4353,N4354);
nor U1593 (N4408,N4355,N4356);
nor U1594 (N4411,N4357,N4358);
nor U1595 (N4414,N4359,N4360);
nor U1596 (N4417,N4361,N4362);
nor U1597 (N4420,N4363,N4364);
nor U1598 (N4423,N4365,N861);
nor U1599 (N4427,N4320,N4368);
nor U1600 (N4428,N4368,N909);
nor U1601 (N4429,N4211,N4368);
nor U1602 (N4432,N4372,N4373);
nor U1603 (N4435,N4377,N4374);
nor U1604 (N4439,N4332,N4380);
nor U1605 (N4440,N4380,N4329);
nor U1606 (N4441,N4384,N4385);
nor U1607 (N4444,N4386,N1104);
nor U1608 (N4448,N4341,N4389);
nor U1609 (N4449,N4389,N1152);
nor U1610 (N4450,N4232,N4389);
nor U1611 (N4453,N4393,N4394);
nor U1612 (N4456,N4398,N4395);
nor U1613 (N4460,N1296,N4401);
nor U1614 (N4461,N4401,N4350);
nor U1615 (N4462,N4405,N573);
nor U1616 (N4466,N4408,N621);
nor U1617 (N4470,N4411,N669);
nor U1618 (N4474,N4414,N717);
nor U1619 (N4478,N4417,N765);
nor U1620 (N4482,N4420,N813);
nor U1621 (N4486,N4365,N4423);
nor U1622 (N4487,N4423,N861);
nor U1623 (N4488,N4260,N4423);
nor U1624 (N4491,N4427,N4428);
nor U1625 (N4494,N4432,N4429);
nor U1626 (N4498,N4377,N4435);
nor U1627 (N4499,N4435,N4374);
nor U1628 (N4500,N4439,N4440);
nor U1629 (N4503,N4441,N1056);
nor U1630 (N4507,N4386,N4444);
nor U1631 (N4508,N4444,N1104);
nor U1632 (N4509,N4281,N4444);
nor U1633 (N4512,N4448,N4449);
nor U1634 (N4515,N4453,N4450);
nor U1635 (N4519,N4398,N4456);
nor U1636 (N4520,N4456,N4395);
nor U1637 (N4521,N4460,N4461);
nor U1638 (N4524,N4405,N4462);
nor U1639 (N4525,N4462,N573);
nor U1640 (N4526,N4294,N4462);
nor U1641 (N4529,N4408,N4466);
nor U1642 (N4530,N4466,N621);
nor U1643 (N4531,N4298,N4466);
nor U1644 (N4534,N4411,N4470);
nor U1645 (N4535,N4470,N669);
nor U1646 (N4536,N4302,N4470);
nor U1647 (N4539,N4414,N4474);
nor U1648 (N4540,N4474,N717);
nor U1649 (N4541,N4306,N4474);
nor U1650 (N4544,N4417,N4478);
nor U1651 (N4545,N4478,N765);
nor U1652 (N4546,N4310,N4478);
nor U1653 (N4549,N4420,N4482);
nor U1654 (N4550,N4482,N813);
nor U1655 (N4551,N4314,N4482);
nor U1656 (N4554,N4486,N4487);
nor U1657 (N4557,N4491,N4488);
nor U1658 (N4561,N4432,N4494);
nor U1659 (N4562,N4494,N4429);
nor U1660 (N4563,N4498,N4499);
nor U1661 (N4566,N4500,N1008);
nor U1662 (N4570,N4441,N4503);
nor U1663 (N4571,N4503,N1056);
nor U1664 (N4572,N4335,N4503);
nor U1665 (N4575,N4507,N4508);
nor U1666 (N4578,N4512,N4509);
nor U1667 (N4582,N4453,N4515);
nor U1668 (N4583,N4515,N4450);
nor U1669 (N4584,N4519,N4520);
nor U1670 (N4587,N4521,N1251);
nor U1671 (N4591,N4524,N4525);
nor U1672 (N4592,N4529,N4530);
nor U1673 (N4595,N4534,N4535);
nor U1674 (N4598,N4539,N4540);
nor U1675 (N4601,N4544,N4545);
nor U1676 (N4604,N4549,N4550);
nor U1677 (N4607,N4554,N4551);
nor U1678 (N4611,N4491,N4557);
nor U1679 (N4612,N4557,N4488);
nor U1680 (N4613,N4561,N4562);
nor U1681 (N4616,N4563,N960);
nor U1682 (N4620,N4500,N4566);
nor U1683 (N4621,N4566,N1008);
nor U1684 (N4622,N4380,N4566);
nor U1685 (N4625,N4570,N4571);
nor U1686 (N4628,N4575,N4572);
nor U1687 (N4632,N4512,N4578);
nor U1688 (N4633,N4578,N4509);
nor U1689 (N4634,N4582,N4583);
nor U1690 (N4637,N4584,N1203);
nor U1691 (N4641,N4521,N4587);
nor U1692 (N4642,N4587,N1251);
nor U1693 (N4643,N4401,N4587);
nor U1694 (N4646,N4592,N4526);
nor U1695 (N4650,N4595,N4531);
nor U1696 (N4654,N4598,N4536);
nor U1697 (N4658,N4601,N4541);
nor U1698 (N4662,N4604,N4546);
nor U1699 (N4666,N4554,N4607);
nor U1700 (N4667,N4607,N4551);
nor U1701 (N4668,N4611,N4612);
nor U1702 (N4671,N4613,N912);
nor U1703 (N4675,N4563,N4616);
nor U1704 (N4676,N4616,N960);
nor U1705 (N4677,N4435,N4616);
nor U1706 (N4680,N4620,N4621);
nor U1707 (N4683,N4625,N4622);
nor U1708 (N4687,N4575,N4628);
nor U1709 (N4688,N4628,N4572);
nor U1710 (N4689,N4632,N4633);
nor U1711 (N4692,N4634,N1155);
nor U1712 (N4696,N4584,N4637);
nor U1713 (N4697,N4637,N1203);
nor U1714 (N4698,N4456,N4637);
nor U1715 (N4701,N4641,N4642);
nor U1716 (N4704,N1299,N4643);
nor U1717 (N4708,N4592,N4646);
nor U1718 (N4709,N4646,N4526);
nor U1719 (N4710,N4595,N4650);
nor U1720 (N4711,N4650,N4531);
nor U1721 (N4712,N4598,N4654);
nor U1722 (N4713,N4654,N4536);
nor U1723 (N4714,N4601,N4658);
nor U1724 (N4715,N4658,N4541);
nor U1725 (N4716,N4604,N4662);
nor U1726 (N4717,N4662,N4546);
nor U1727 (N4718,N4666,N4667);
nor U1728 (N4721,N4668,N864);
nor U1729 (N4725,N4613,N4671);
nor U1730 (N4726,N4671,N912);
nor U1731 (N4727,N4494,N4671);
nor U1732 (N4730,N4675,N4676);
nor U1733 (N4733,N4680,N4677);
nor U1734 (N4737,N4625,N4683);
nor U1735 (N4738,N4683,N4622);
nor U1736 (N4739,N4687,N4688);
nor U1737 (N4742,N4689,N1107);
nor U1738 (N4746,N4634,N4692);
nor U1739 (N4747,N4692,N1155);
nor U1740 (N4748,N4515,N4692);
nor U1741 (N4751,N4696,N4697);
nor U1742 (N4754,N4701,N4698);
nor U1743 (N4758,N1299,N4704);
nor U1744 (N4759,N4704,N4643);
nor U1745 (N4760,N4708,N4709);
nor U1746 (N4763,N4710,N4711);
nor U1747 (N4766,N4712,N4713);
nor U1748 (N4769,N4714,N4715);
nor U1749 (N4772,N4716,N4717);
nor U1750 (N4775,N4718,N816);
nor U1751 (N4779,N4668,N4721);
nor U1752 (N4780,N4721,N864);
nor U1753 (N4781,N4557,N4721);
nor U1754 (N4784,N4725,N4726);
nor U1755 (N4787,N4730,N4727);
nor U1756 (N4791,N4680,N4733);
nor U1757 (N4792,N4733,N4677);
nor U1758 (N4793,N4737,N4738);
nor U1759 (N4796,N4739,N1059);
nor U1760 (N4800,N4689,N4742);
nor U1761 (N4801,N4742,N1107);
nor U1762 (N4802,N4578,N4742);
nor U1763 (N4805,N4746,N4747);
nor U1764 (N4808,N4751,N4748);
nor U1765 (N4812,N4701,N4754);
nor U1766 (N4813,N4754,N4698);
nor U1767 (N4814,N4758,N4759);
nor U1768 (N4817,N4760,N576);
nor U1769 (N4821,N4763,N624);
nor U1770 (N4825,N4766,N672);
nor U1771 (N4829,N4769,N720);
nor U1772 (N4833,N4772,N768);
nor U1773 (N4837,N4718,N4775);
nor U1774 (N4838,N4775,N816);
nor U1775 (N4839,N4607,N4775);
nor U1776 (N4842,N4779,N4780);
nor U1777 (N4845,N4784,N4781);
nor U1778 (N4849,N4730,N4787);
nor U1779 (N4850,N4787,N4727);
nor U1780 (N4851,N4791,N4792);
nor U1781 (N4854,N4793,N1011);
nor U1782 (N4858,N4739,N4796);
nor U1783 (N4859,N4796,N1059);
nor U1784 (N4860,N4628,N4796);
nor U1785 (N4863,N4800,N4801);
nor U1786 (N4866,N4805,N4802);
nor U1787 (N4870,N4751,N4808);
nor U1788 (N4871,N4808,N4748);
nor U1789 (N4872,N4812,N4813);
nor U1790 (N4875,N4814,N1254);
nor U1791 (N4879,N4760,N4817);
nor U1792 (N4880,N4817,N576);
nor U1793 (N4881,N4646,N4817);
nor U1794 (N4884,N4763,N4821);
nor U1795 (N4885,N4821,N624);
nor U1796 (N4886,N4650,N4821);
nor U1797 (N4889,N4766,N4825);
nor U1798 (N4890,N4825,N672);
nor U1799 (N4891,N4654,N4825);
nor U1800 (N4894,N4769,N4829);
nor U1801 (N4895,N4829,N720);
nor U1802 (N4896,N4658,N4829);
nor U1803 (N4899,N4772,N4833);
nor U1804 (N4900,N4833,N768);
nor U1805 (N4901,N4662,N4833);
nor U1806 (N4904,N4837,N4838);
nor U1807 (N4907,N4842,N4839);
nor U1808 (N4911,N4784,N4845);
nor U1809 (N4912,N4845,N4781);
nor U1810 (N4913,N4849,N4850);
nor U1811 (N4916,N4851,N963);
nor U1812 (N4920,N4793,N4854);
nor U1813 (N4921,N4854,N1011);
nor U1814 (N4922,N4683,N4854);
nor U1815 (N4925,N4858,N4859);
nor U1816 (N4928,N4863,N4860);
nor U1817 (N4932,N4805,N4866);
nor U1818 (N4933,N4866,N4802);
nor U1819 (N4934,N4870,N4871);
nor U1820 (N4937,N4872,N1206);
nor U1821 (N4941,N4814,N4875);
nor U1822 (N4942,N4875,N1254);
nor U1823 (N4943,N4704,N4875);
nor U1824 (N4946,N4879,N4880);
nor U1825 (N4947,N4884,N4885);
nor U1826 (N4950,N4889,N4890);
nor U1827 (N4953,N4894,N4895);
nor U1828 (N4956,N4899,N4900);
nor U1829 (N4959,N4904,N4901);
nor U1830 (N4963,N4842,N4907);
nor U1831 (N4964,N4907,N4839);
nor U1832 (N4965,N4911,N4912);
nor U1833 (N4968,N4913,N915);
nor U1834 (N4972,N4851,N4916);
nor U1835 (N4973,N4916,N963);
nor U1836 (N4974,N4733,N4916);
nor U1837 (N4977,N4920,N4921);
nor U1838 (N4980,N4925,N4922);
nor U1839 (N4984,N4863,N4928);
nor U1840 (N4985,N4928,N4860);
nor U1841 (N4986,N4932,N4933);
nor U1842 (N4989,N4934,N1158);
nor U1843 (N4993,N4872,N4937);
nor U1844 (N4994,N4937,N1206);
nor U1845 (N4995,N4754,N4937);
nor U1846 (N4998,N4941,N4942);
nor U1847 (N5001,N1302,N4943);
nor U1848 (N5005,N4947,N4881);
nor U1849 (N5009,N4950,N4886);
nor U1850 (N5013,N4953,N4891);
nor U1851 (N5017,N4956,N4896);
nor U1852 (N5021,N4904,N4959);
nor U1853 (N5022,N4959,N4901);
nor U1854 (N5023,N4963,N4964);
nor U1855 (N5026,N4965,N867);
nor U1856 (N5030,N4913,N4968);
nor U1857 (N5031,N4968,N915);
nor U1858 (N5032,N4787,N4968);
nor U1859 (N5035,N4972,N4973);
nor U1860 (N5038,N4977,N4974);
nor U1861 (N5042,N4925,N4980);
nor U1862 (N5043,N4980,N4922);
nor U1863 (N5044,N4984,N4985);
nor U1864 (N5047,N4986,N1110);
nor U1865 (N5051,N4934,N4989);
nor U1866 (N5052,N4989,N1158);
nor U1867 (N5053,N4808,N4989);
nor U1868 (N5056,N4993,N4994);
nor U1869 (N5059,N4998,N4995);
nor U1870 (N5063,N1302,N5001);
nor U1871 (N5064,N5001,N4943);
nor U1872 (N5065,N4947,N5005);
nor U1873 (N5066,N5005,N4881);
nor U1874 (N5067,N4950,N5009);
nor U1875 (N5068,N5009,N4886);
nor U1876 (N5069,N4953,N5013);
nor U1877 (N5070,N5013,N4891);
nor U1878 (N5071,N4956,N5017);
nor U1879 (N5072,N5017,N4896);
nor U1880 (N5073,N5021,N5022);
nor U1881 (N5076,N5023,N819);
nor U1882 (N5080,N4965,N5026);
nor U1883 (N5081,N5026,N867);
nor U1884 (N5082,N4845,N5026);
nor U1885 (N5085,N5030,N5031);
nor U1886 (N5088,N5035,N5032);
nor U1887 (N5092,N4977,N5038);
nor U1888 (N5093,N5038,N4974);
nor U1889 (N5094,N5042,N5043);
nor U1890 (N5097,N5044,N1062);
nor U1891 (N5101,N4986,N5047);
nor U1892 (N5102,N5047,N1110);
nor U1893 (N5103,N4866,N5047);
nor U1894 (N5106,N5051,N5052);
nor U1895 (N5109,N5056,N5053);
nor U1896 (N5113,N4998,N5059);
nor U1897 (N5114,N5059,N4995);
nor U1898 (N5115,N5063,N5064);
nor U1899 (N5118,N5065,N5066);
nor U1900 (N5121,N5067,N5068);
nor U1901 (N5124,N5069,N5070);
nor U1902 (N5127,N5071,N5072);
nor U1903 (N5130,N5073,N771);
nor U1904 (N5134,N5023,N5076);
nor U1905 (N5135,N5076,N819);
nor U1906 (N5136,N4907,N5076);
nor U1907 (N5139,N5080,N5081);
nor U1908 (N5142,N5085,N5082);
nor U1909 (N5146,N5035,N5088);
nor U1910 (N5147,N5088,N5032);
nor U1911 (N5148,N5092,N5093);
nor U1912 (N5151,N5094,N1014);
nor U1913 (N5155,N5044,N5097);
nor U1914 (N5156,N5097,N1062);
nor U1915 (N5157,N4928,N5097);
nor U1916 (N5160,N5101,N5102);
nor U1917 (N5163,N5106,N5103);
nor U1918 (N5167,N5056,N5109);
nor U1919 (N5168,N5109,N5053);
nor U1920 (N5169,N5113,N5114);
nor U1921 (N5172,N5115,N1257);
nor U1922 (N5176,N5118,N579);
nor U1923 (N5180,N5121,N627);
nor U1924 (N5184,N5124,N675);
nor U1925 (N5188,N5127,N723);
nor U1926 (N5192,N5073,N5130);
nor U1927 (N5193,N5130,N771);
nor U1928 (N5194,N4959,N5130);
nor U1929 (N5197,N5134,N5135);
nor U1930 (N5200,N5139,N5136);
nor U1931 (N5204,N5085,N5142);
nor U1932 (N5205,N5142,N5082);
nor U1933 (N5206,N5146,N5147);
nor U1934 (N5209,N5148,N966);
nor U1935 (N5213,N5094,N5151);
nor U1936 (N5214,N5151,N1014);
nor U1937 (N5215,N4980,N5151);
nor U1938 (N5218,N5155,N5156);
nor U1939 (N5221,N5160,N5157);
nor U1940 (N5225,N5106,N5163);
nor U1941 (N5226,N5163,N5103);
nor U1942 (N5227,N5167,N5168);
nor U1943 (N5230,N5169,N1209);
nor U1944 (N5234,N5115,N5172);
nor U1945 (N5235,N5172,N1257);
nor U1946 (N5236,N5001,N5172);
nor U1947 (N5239,N5118,N5176);
nor U1948 (N5240,N5176,N579);
nor U1949 (N5241,N5005,N5176);
nor U1950 (N5244,N5121,N5180);
nor U1951 (N5245,N5180,N627);
nor U1952 (N5246,N5009,N5180);
nor U1953 (N5249,N5124,N5184);
nor U1954 (N5250,N5184,N675);
nor U1955 (N5251,N5013,N5184);
nor U1956 (N5254,N5127,N5188);
nor U1957 (N5255,N5188,N723);
nor U1958 (N5256,N5017,N5188);
nor U1959 (N5259,N5192,N5193);
nor U1960 (N5262,N5197,N5194);
nor U1961 (N5266,N5139,N5200);
nor U1962 (N5267,N5200,N5136);
nor U1963 (N5268,N5204,N5205);
nor U1964 (N5271,N5206,N918);
nor U1965 (N5275,N5148,N5209);
nor U1966 (N5276,N5209,N966);
nor U1967 (N5277,N5038,N5209);
nor U1968 (N5280,N5213,N5214);
nor U1969 (N5283,N5218,N5215);
nor U1970 (N5287,N5160,N5221);
nor U1971 (N5288,N5221,N5157);
nor U1972 (N5289,N5225,N5226);
nor U1973 (N5292,N5227,N1161);
nor U1974 (N5296,N5169,N5230);
nor U1975 (N5297,N5230,N1209);
nor U1976 (N5298,N5059,N5230);
nor U1977 (N5301,N5234,N5235);
nor U1978 (N5304,N1305,N5236);
nor U1979 (N5308,N5239,N5240);
nor U1980 (N5309,N5244,N5245);
nor U1981 (N5312,N5249,N5250);
nor U1982 (N5315,N5254,N5255);
nor U1983 (N5318,N5259,N5256);
nor U1984 (N5322,N5197,N5262);
nor U1985 (N5323,N5262,N5194);
nor U1986 (N5324,N5266,N5267);
nor U1987 (N5327,N5268,N870);
nor U1988 (N5331,N5206,N5271);
nor U1989 (N5332,N5271,N918);
nor U1990 (N5333,N5088,N5271);
nor U1991 (N5336,N5275,N5276);
nor U1992 (N5339,N5280,N5277);
nor U1993 (N5343,N5218,N5283);
nor U1994 (N5344,N5283,N5215);
nor U1995 (N5345,N5287,N5288);
nor U1996 (N5348,N5289,N1113);
nor U1997 (N5352,N5227,N5292);
nor U1998 (N5353,N5292,N1161);
nor U1999 (N5354,N5109,N5292);
nor U2000 (N5357,N5296,N5297);
nor U2001 (N5360,N5301,N5298);
nor U2002 (N5364,N1305,N5304);
nor U2003 (N5365,N5304,N5236);
nor U2004 (N5366,N5309,N5241);
nor U2005 (N5370,N5312,N5246);
nor U2006 (N5374,N5315,N5251);
nor U2007 (N5378,N5259,N5318);
nor U2008 (N5379,N5318,N5256);
nor U2009 (N5380,N5322,N5323);
nor U2010 (N5383,N5324,N822);
nor U2011 (N5387,N5268,N5327);
nor U2012 (N5388,N5327,N870);
nor U2013 (N5389,N5142,N5327);
nor U2014 (N5392,N5331,N5332);
nor U2015 (N5395,N5336,N5333);
nor U2016 (N5399,N5280,N5339);
nor U2017 (N5400,N5339,N5277);
nor U2018 (N5401,N5343,N5344);
nor U2019 (N5404,N5345,N1065);
nor U2020 (N5408,N5289,N5348);
nor U2021 (N5409,N5348,N1113);
nor U2022 (N5410,N5163,N5348);
nor U2023 (N5413,N5352,N5353);
nor U2024 (N5416,N5357,N5354);
nor U2025 (N5420,N5301,N5360);
nor U2026 (N5421,N5360,N5298);
nor U2027 (N5422,N5364,N5365);
nor U2028 (N5425,N5309,N5366);
nor U2029 (N5426,N5366,N5241);
nor U2030 (N5427,N5312,N5370);
nor U2031 (N5428,N5370,N5246);
nor U2032 (N5429,N5315,N5374);
nor U2033 (N5430,N5374,N5251);
nor U2034 (N5431,N5378,N5379);
nor U2035 (N5434,N5380,N774);
nor U2036 (N5438,N5324,N5383);
nor U2037 (N5439,N5383,N822);
nor U2038 (N5440,N5200,N5383);
nor U2039 (N5443,N5387,N5388);
nor U2040 (N5446,N5392,N5389);
nor U2041 (N5450,N5336,N5395);
nor U2042 (N5451,N5395,N5333);
nor U2043 (N5452,N5399,N5400);
nor U2044 (N5455,N5401,N1017);
nor U2045 (N5459,N5345,N5404);
nor U2046 (N5460,N5404,N1065);
nor U2047 (N5461,N5221,N5404);
nor U2048 (N5464,N5408,N5409);
nor U2049 (N5467,N5413,N5410);
nor U2050 (N5471,N5357,N5416);
nor U2051 (N5472,N5416,N5354);
nor U2052 (N5473,N5420,N5421);
nor U2053 (N5476,N5422,N1260);
nor U2054 (N5480,N5425,N5426);
nor U2055 (N5483,N5427,N5428);
nor U2056 (N5486,N5429,N5430);
nor U2057 (N5489,N5431,N726);
nor U2058 (N5493,N5380,N5434);
nor U2059 (N5494,N5434,N774);
nor U2060 (N5495,N5262,N5434);
nor U2061 (N5498,N5438,N5439);
nor U2062 (N5501,N5443,N5440);
nor U2063 (N5505,N5392,N5446);
nor U2064 (N5506,N5446,N5389);
nor U2065 (N5507,N5450,N5451);
nor U2066 (N5510,N5452,N969);
nor U2067 (N5514,N5401,N5455);
nor U2068 (N5515,N5455,N1017);
nor U2069 (N5516,N5283,N5455);
nor U2070 (N5519,N5459,N5460);
nor U2071 (N5522,N5464,N5461);
nor U2072 (N5526,N5413,N5467);
nor U2073 (N5527,N5467,N5410);
nor U2074 (N5528,N5471,N5472);
nor U2075 (N5531,N5473,N1212);
nor U2076 (N5535,N5422,N5476);
nor U2077 (N5536,N5476,N1260);
nor U2078 (N5537,N5304,N5476);
nor U2079 (N5540,N5480,N582);
nor U2080 (N5544,N5483,N630);
nor U2081 (N5548,N5486,N678);
nor U2082 (N5552,N5431,N5489);
nor U2083 (N5553,N5489,N726);
nor U2084 (N5554,N5318,N5489);
nor U2085 (N5557,N5493,N5494);
nor U2086 (N5560,N5498,N5495);
nor U2087 (N5564,N5443,N5501);
nor U2088 (N5565,N5501,N5440);
nor U2089 (N5566,N5505,N5506);
nor U2090 (N5569,N5507,N921);
nor U2091 (N5573,N5452,N5510);
nor U2092 (N5574,N5510,N969);
nor U2093 (N5575,N5339,N5510);
nor U2094 (N5578,N5514,N5515);
nor U2095 (N5581,N5519,N5516);
nor U2096 (N5585,N5464,N5522);
nor U2097 (N5586,N5522,N5461);
nor U2098 (N5587,N5526,N5527);
nor U2099 (N5590,N5528,N1164);
nor U2100 (N5594,N5473,N5531);
nor U2101 (N5595,N5531,N1212);
nor U2102 (N5596,N5360,N5531);
nor U2103 (N5599,N5535,N5536);
nor U2104 (N5602,N1308,N5537);
nor U2105 (N5606,N5480,N5540);
nor U2106 (N5607,N5540,N582);
nor U2107 (N5608,N5366,N5540);
nor U2108 (N5611,N5483,N5544);
nor U2109 (N5612,N5544,N630);
nor U2110 (N5613,N5370,N5544);
nor U2111 (N5616,N5486,N5548);
nor U2112 (N5617,N5548,N678);
nor U2113 (N5618,N5374,N5548);
nor U2114 (N5621,N5552,N5553);
nor U2115 (N5624,N5557,N5554);
nor U2116 (N5628,N5498,N5560);
nor U2117 (N5629,N5560,N5495);
nor U2118 (N5630,N5564,N5565);
nor U2119 (N5633,N5566,N873);
nor U2120 (N5637,N5507,N5569);
nor U2121 (N5638,N5569,N921);
nor U2122 (N5639,N5395,N5569);
nor U2123 (N5642,N5573,N5574);
nor U2124 (N5645,N5578,N5575);
nor U2125 (N5649,N5519,N5581);
nor U2126 (N5650,N5581,N5516);
nor U2127 (N5651,N5585,N5586);
nor U2128 (N5654,N5587,N1116);
nor U2129 (N5658,N5528,N5590);
nor U2130 (N5659,N5590,N1164);
nor U2131 (N5660,N5416,N5590);
nor U2132 (N5663,N5594,N5595);
nor U2133 (N5666,N5599,N5596);
nor U2134 (N5670,N1308,N5602);
nor U2135 (N5671,N5602,N5537);
nor U2136 (N5672,N5606,N5607);
nor U2137 (N5673,N5611,N5612);
nor U2138 (N5676,N5616,N5617);
nor U2139 (N5679,N5621,N5618);
nor U2140 (N5683,N5557,N5624);
nor U2141 (N5684,N5624,N5554);
nor U2142 (N5685,N5628,N5629);
nor U2143 (N5688,N5630,N825);
nor U2144 (N5692,N5566,N5633);
nor U2145 (N5693,N5633,N873);
nor U2146 (N5694,N5446,N5633);
nor U2147 (N5697,N5637,N5638);
nor U2148 (N5700,N5642,N5639);
nor U2149 (N5704,N5578,N5645);
nor U2150 (N5705,N5645,N5575);
nor U2151 (N5706,N5649,N5650);
nor U2152 (N5709,N5651,N1068);
nor U2153 (N5713,N5587,N5654);
nor U2154 (N5714,N5654,N1116);
nor U2155 (N5715,N5467,N5654);
nor U2156 (N5718,N5658,N5659);
nor U2157 (N5721,N5663,N5660);
nor U2158 (N5725,N5599,N5666);
nor U2159 (N5726,N5666,N5596);
nor U2160 (N5727,N5670,N5671);
nor U2161 (N5730,N5673,N5608);
nor U2162 (N5734,N5676,N5613);
nor U2163 (N5738,N5621,N5679);
nor U2164 (N5739,N5679,N5618);
nor U2165 (N5740,N5683,N5684);
nor U2166 (N5743,N5685,N777);
nor U2167 (N5747,N5630,N5688);
nor U2168 (N5748,N5688,N825);
nor U2169 (N5749,N5501,N5688);
nor U2170 (N5752,N5692,N5693);
nor U2171 (N5755,N5697,N5694);
nor U2172 (N5759,N5642,N5700);
nor U2173 (N5760,N5700,N5639);
nor U2174 (N5761,N5704,N5705);
nor U2175 (N5764,N5706,N1020);
nor U2176 (N5768,N5651,N5709);
nor U2177 (N5769,N5709,N1068);
nor U2178 (N5770,N5522,N5709);
nor U2179 (N5773,N5713,N5714);
nor U2180 (N5776,N5718,N5715);
nor U2181 (N5780,N5663,N5721);
nor U2182 (N5781,N5721,N5660);
nor U2183 (N5782,N5725,N5726);
nor U2184 (N5785,N5673,N5730);
nor U2185 (N5786,N5730,N5608);
nor U2186 (N5787,N5676,N5734);
nor U2187 (N5788,N5734,N5613);
nor U2188 (N5789,N5738,N5739);
nor U2189 (N5792,N5740,N729);
nor U2190 (N5796,N5685,N5743);
nor U2191 (N5797,N5743,N777);
nor U2192 (N5798,N5560,N5743);
nor U2193 (N5801,N5747,N5748);
nor U2194 (N5804,N5752,N5749);
nor U2195 (N5808,N5697,N5755);
nor U2196 (N5809,N5755,N5694);
nor U2197 (N5810,N5759,N5760);
nor U2198 (N5813,N5761,N972);
nor U2199 (N5817,N5706,N5764);
nor U2200 (N5818,N5764,N1020);
nor U2201 (N5819,N5581,N5764);
nor U2202 (N5822,N5768,N5769);
nor U2203 (N5825,N5773,N5770);
nor U2204 (N5829,N5718,N5776);
nor U2205 (N5830,N5776,N5715);
nor U2206 (N5831,N5780,N5781);
nor U2207 (N5834,N5785,N5786);
nor U2208 (N5837,N5787,N5788);
nor U2209 (N5840,N5789,N681);
nor U2210 (N5844,N5740,N5792);
nor U2211 (N5845,N5792,N729);
nor U2212 (N5846,N5624,N5792);
nor U2213 (N5849,N5796,N5797);
nor U2214 (N5852,N5801,N5798);
nor U2215 (N5856,N5752,N5804);
nor U2216 (N5857,N5804,N5749);
nor U2217 (N5858,N5808,N5809);
nor U2218 (N5861,N5810,N924);
nor U2219 (N5865,N5761,N5813);
nor U2220 (N5866,N5813,N972);
nor U2221 (N5867,N5645,N5813);
nor U2222 (N5870,N5817,N5818);
nor U2223 (N5873,N5822,N5819);
nor U2224 (N5877,N5773,N5825);
nor U2225 (N5878,N5825,N5770);
nor U2226 (N5879,N5829,N5830);
nor U2227 (N5882,N5834,N585);
nor U2228 (N5886,N5837,N633);
nor U2229 (N5890,N5789,N5840);
nor U2230 (N5891,N5840,N681);
nor U2231 (N5892,N5679,N5840);
nor U2232 (N5895,N5844,N5845);
nor U2233 (N5898,N5849,N5846);
nor U2234 (N5902,N5801,N5852);
nor U2235 (N5903,N5852,N5798);
nor U2236 (N5904,N5856,N5857);
nor U2237 (N5907,N5858,N876);
nor U2238 (N5911,N5810,N5861);
nor U2239 (N5912,N5861,N924);
nor U2240 (N5913,N5700,N5861);
nor U2241 (N5916,N5865,N5866);
nor U2242 (N5919,N5870,N5867);
nor U2243 (N5923,N5822,N5873);
nor U2244 (N5924,N5873,N5819);
nor U2245 (N5925,N5877,N5878);
nor U2246 (N5928,N5834,N5882);
nor U2247 (N5929,N5882,N585);
nor U2248 (N5930,N5730,N5882);
nor U2249 (N5933,N5837,N5886);
nor U2250 (N5934,N5886,N633);
nor U2251 (N5935,N5734,N5886);
nor U2252 (N5938,N5890,N5891);
nor U2253 (N5941,N5895,N5892);
nor U2254 (N5945,N5849,N5898);
nor U2255 (N5946,N5898,N5846);
nor U2256 (N5947,N5902,N5903);
nor U2257 (N5950,N5904,N828);
nor U2258 (N5954,N5858,N5907);
nor U2259 (N5955,N5907,N876);
nor U2260 (N5956,N5755,N5907);
nor U2261 (N5959,N5911,N5912);
nor U2262 (N5962,N5916,N5913);
nor U2263 (N5966,N5870,N5919);
nor U2264 (N5967,N5919,N5867);
nor U2265 (N5968,N5923,N5924);
nor U2266 (N5971,N5928,N5929);
nor U2267 (N5972,N5933,N5934);
nor U2268 (N5975,N5938,N5935);
nor U2269 (N5979,N5895,N5941);
nor U2270 (N5980,N5941,N5892);
nor U2271 (N5981,N5945,N5946);
nor U2272 (N5984,N5947,N780);
nor U2273 (N5988,N5904,N5950);
nor U2274 (N5989,N5950,N828);
nor U2275 (N5990,N5804,N5950);
nor U2276 (N5993,N5954,N5955);
nor U2277 (N5996,N5959,N5956);
nor U2278 (N6000,N5916,N5962);
nor U2279 (N6001,N5962,N5913);
nor U2280 (N6002,N5966,N5967);
nor U2281 (N6005,N5972,N5930);
nor U2282 (N6009,N5938,N5975);
nor U2283 (N6010,N5975,N5935);
nor U2284 (N6011,N5979,N5980);
nor U2285 (N6014,N5981,N732);
nor U2286 (N6018,N5947,N5984);
nor U2287 (N6019,N5984,N780);
nor U2288 (N6020,N5852,N5984);
nor U2289 (N6023,N5988,N5989);
nor U2290 (N6026,N5993,N5990);
nor U2291 (N6030,N5959,N5996);
nor U2292 (N6031,N5996,N5956);
nor U2293 (N6032,N6000,N6001);
nor U2294 (N6035,N5972,N6005);
nor U2295 (N6036,N6005,N5930);
nor U2296 (N6037,N6009,N6010);
nor U2297 (N6040,N6011,N684);
nor U2298 (N6044,N5981,N6014);
nor U2299 (N6045,N6014,N732);
nor U2300 (N6046,N5898,N6014);
nor U2301 (N6049,N6018,N6019);
nor U2302 (N6052,N6023,N6020);
nor U2303 (N6056,N5993,N6026);
nor U2304 (N6057,N6026,N5990);
nor U2305 (N6058,N6030,N6031);
nor U2306 (N6061,N6035,N6036);
nor U2307 (N6064,N6037,N636);
nor U2308 (N6068,N6011,N6040);
nor U2309 (N6069,N6040,N684);
nor U2310 (N6070,N5941,N6040);
nor U2311 (N6073,N6044,N6045);
nor U2312 (N6076,N6049,N6046);
nor U2313 (N6080,N6023,N6052);
nor U2314 (N6081,N6052,N6020);
nor U2315 (N6082,N6056,N6057);
nor U2316 (N6085,N6061,N588);
nor U2317 (N6089,N6037,N6064);
nor U2318 (N6090,N6064,N636);
nor U2319 (N6091,N5975,N6064);
nor U2320 (N6094,N6068,N6069);
nor U2321 (N6097,N6073,N6070);
nor U2322 (N6101,N6049,N6076);
nor U2323 (N6102,N6076,N6046);
nor U2324 (N6103,N6080,N6081);
nor U2325 (N6106,N6061,N6085);
nor U2326 (N6107,N6085,N588);
nor U2327 (N6108,N6005,N6085);
nor U2328 (N6111,N6089,N6090);
nor U2329 (N6114,N6094,N6091);
nor U2330 (N6118,N6073,N6097);
nor U2331 (N6119,N6097,N6070);
nor U2332 (N6120,N6101,N6102);
nor U2333 (N6123,N6106,N6107);
nor U2334 (N6124,N6111,N6108);
nor U2335 (N6128,N6094,N6114);
nor U2336 (N6129,N6114,N6091);
nor U2337 (N6130,N6118,N6119);
nor U2338 (N6133,N6111,N6124);
nor U2339 (N6134,N6124,N6108);
nor U2340 (N6135,N6128,N6129);
nor U2341 (N6138,N6133,N6134);
not U2342 (N6141,N6138);
nor U2343 (N6145,N6138,N6141);
not U2344 (N6146,N6141);
nor U2345 (N6147,N6124,N6141);
nor U2346 (N6150,N6145,N6146);
nor U2347 (N6151,N6135,N6147);
nor U2348 (N6155,N6135,N6151);
nor U2349 (N6156,N6151,N6147);
nor U2350 (N6157,N6114,N6151);
nor U2351 (N6160,N6155,N6156);
nor U2352 (N6161,N6130,N6157);
nor U2353 (N6165,N6130,N6161);
nor U2354 (N6166,N6161,N6157);
nor U2355 (N6167,N6097,N6161);
nor U2356 (N6170,N6165,N6166);
nor U2357 (N6171,N6120,N6167);
nor U2358 (N6175,N6120,N6171);
nor U2359 (N6176,N6171,N6167);
nor U2360 (N6177,N6076,N6171);
nor U2361 (N6180,N6175,N6176);
nor U2362 (N6181,N6103,N6177);
nor U2363 (N6185,N6103,N6181);
nor U2364 (N6186,N6181,N6177);
nor U2365 (N6187,N6052,N6181);
nor U2366 (N6190,N6185,N6186);
nor U2367 (N6191,N6082,N6187);
nor U2368 (N6195,N6082,N6191);
nor U2369 (N6196,N6191,N6187);
nor U2370 (N6197,N6026,N6191);
nor U2371 (N6200,N6195,N6196);
nor U2372 (N6201,N6058,N6197);
nor U2373 (N6205,N6058,N6201);
nor U2374 (N6206,N6201,N6197);
nor U2375 (N6207,N5996,N6201);
nor U2376 (N6210,N6205,N6206);
nor U2377 (N6211,N6032,N6207);
nor U2378 (N6215,N6032,N6211);
nor U2379 (N6216,N6211,N6207);
nor U2380 (N6217,N5962,N6211);
nor U2381 (N6220,N6215,N6216);
nor U2382 (N6221,N6002,N6217);
nor U2383 (N6225,N6002,N6221);
nor U2384 (N6226,N6221,N6217);
nor U2385 (N6227,N5919,N6221);
nor U2386 (N6230,N6225,N6226);
nor U2387 (N6231,N5968,N6227);
nor U2388 (N6235,N5968,N6231);
nor U2389 (N6236,N6231,N6227);
nor U2390 (N6237,N5873,N6231);
nor U2391 (N6240,N6235,N6236);
nor U2392 (N6241,N5925,N6237);
nor U2393 (N6245,N5925,N6241);
nor U2394 (N6246,N6241,N6237);
nor U2395 (N6247,N5825,N6241);
nor U2396 (N6250,N6245,N6246);
nor U2397 (N6251,N5879,N6247);
nor U2398 (N6255,N5879,N6251);
nor U2399 (N6256,N6251,N6247);
nor U2400 (N6257,N5776,N6251);
nor U2401 (N6260,N6255,N6256);
nor U2402 (N6261,N5831,N6257);
nor U2403 (N6265,N5831,N6261);
nor U2404 (N6266,N6261,N6257);
nor U2405 (N6267,N5721,N6261);
nor U2406 (N6270,N6265,N6266);
nor U2407 (N6271,N5782,N6267);
nor U2408 (N6275,N5782,N6271);
nor U2409 (N6276,N6271,N6267);
nor U2410 (N6277,N5666,N6271);
nor U2411 (N6280,N6275,N6276);
nor U2412 (N6281,N5727,N6277);
nor U2413 (N6285,N5727,N6281);
nor U2414 (N6286,N6281,N6277);
nor U2415 (N6287,N5602,N6281);
nor U2416 (N6288,N6285,N6286);
endmodule
