module ibex (rst_ni, hart_id_i_31_, hart_id_i_30_, hart_id_i_29_, hart_id_i_28_, hart_id_i_27_, hart_id_i_26_, hart_id_i_25_, hart_id_i_24_, hart_id_i_23_, hart_id_i_22_, hart_id_i_21_, hart_id_i_20_, hart_id_i_19_, hart_id_i_18_, hart_id_i_17_, hart_id_i_16_, hart_id_i_15_, hart_id_i_14_, hart_id_i_13_, hart_id_i_12_, hart_id_i_11_, hart_id_i_10_, hart_id_i_9_, hart_id_i_8_, hart_id_i_7_, hart_id_i_6_, hart_id_i_5_, hart_id_i_4_, hart_id_i_3_, hart_id_i_2_, hart_id_i_1_, hart_id_i_0_, boot_addr_i_31_, boot_addr_i_30_, boot_addr_i_29_, boot_addr_i_28_, boot_addr_i_27_, boot_addr_i_26_, boot_addr_i_25_, boot_addr_i_24_, boot_addr_i_23_, boot_addr_i_22_, boot_addr_i_21_, boot_addr_i_20_, boot_addr_i_19_, boot_addr_i_18_, boot_addr_i_17_, boot_addr_i_16_, boot_addr_i_15_, boot_addr_i_14_, boot_addr_i_13_, boot_addr_i_12_, boot_addr_i_11_, boot_addr_i_10_, boot_addr_i_9_, boot_addr_i_8_, boot_addr_i_7_, boot_addr_i_6_, boot_addr_i_5_, boot_addr_i_4_, boot_addr_i_3_, boot_addr_i_2_, boot_addr_i_1_, boot_addr_i_0_, instr_req_o, instr_gnt_i, instr_rvalid_i, instr_addr_o_31_, instr_addr_o_30_, instr_addr_o_29_, instr_addr_o_28_, instr_addr_o_27_, instr_addr_o_26_, instr_addr_o_25_, instr_addr_o_24_, instr_addr_o_23_, instr_addr_o_22_, instr_addr_o_21_, instr_addr_o_20_, instr_addr_o_19_, instr_addr_o_18_, instr_addr_o_17_, instr_addr_o_16_, instr_addr_o_15_, instr_addr_o_14_, instr_addr_o_13_, instr_addr_o_12_, instr_addr_o_11_, instr_addr_o_10_, instr_addr_o_9_, instr_addr_o_8_, instr_addr_o_7_, instr_addr_o_6_, instr_addr_o_5_, instr_addr_o_4_, instr_addr_o_3_, instr_addr_o_2_, instr_addr_o_1_, instr_addr_o_0_, instr_rdata_i_31_, instr_rdata_i_30_, instr_rdata_i_29_, instr_rdata_i_28_, instr_rdata_i_27_, instr_rdata_i_26_, instr_rdata_i_25_, instr_rdata_i_24_, instr_rdata_i_23_, instr_rdata_i_22_, instr_rdata_i_21_, instr_rdata_i_20_, instr_rdata_i_19_, instr_rdata_i_18_, instr_rdata_i_17_, instr_rdata_i_16_, instr_rdata_i_15_, instr_rdata_i_14_, instr_rdata_i_13_, instr_rdata_i_12_, instr_rdata_i_11_, instr_rdata_i_10_, instr_rdata_i_9_, instr_rdata_i_8_, instr_rdata_i_7_, instr_rdata_i_6_, instr_rdata_i_5_, instr_rdata_i_4_, instr_rdata_i_3_, instr_rdata_i_2_, instr_rdata_i_1_, instr_rdata_i_0_, instr_err_i, data_req_o, data_gnt_i, data_rvalid_i, data_we_o, data_be_o_3_, data_be_o_2_, data_be_o_1_, data_be_o_0_, data_addr_o_31_, data_addr_o_30_, data_addr_o_29_, data_addr_o_28_, data_addr_o_27_, data_addr_o_26_, data_addr_o_25_, data_addr_o_24_, data_addr_o_23_, data_addr_o_22_, data_addr_o_21_, data_addr_o_20_, data_addr_o_19_, data_addr_o_18_, data_addr_o_17_, data_addr_o_16_, data_addr_o_15_, data_addr_o_14_, data_addr_o_13_, data_addr_o_12_, data_addr_o_11_, data_addr_o_10_, data_addr_o_9_, data_addr_o_8_, data_addr_o_7_, data_addr_o_6_, data_addr_o_5_, data_addr_o_4_, data_addr_o_3_, data_addr_o_2_, data_addr_o_1_, data_addr_o_0_, data_wdata_o_31_, data_wdata_o_30_, data_wdata_o_29_, data_wdata_o_28_, data_wdata_o_27_, data_wdata_o_26_, data_wdata_o_25_, data_wdata_o_24_, data_wdata_o_23_, data_wdata_o_22_, data_wdata_o_21_, data_wdata_o_20_, data_wdata_o_19_, data_wdata_o_18_, data_wdata_o_17_, data_wdata_o_16_, data_wdata_o_15_, data_wdata_o_14_, data_wdata_o_13_, data_wdata_o_12_, data_wdata_o_11_, data_wdata_o_10_, data_wdata_o_9_, data_wdata_o_8_, data_wdata_o_7_, data_wdata_o_6_, data_wdata_o_5_, data_wdata_o_4_, data_wdata_o_3_, data_wdata_o_2_, data_wdata_o_1_, data_wdata_o_0_, data_rdata_i_31_, data_rdata_i_30_, data_rdata_i_29_, data_rdata_i_28_, data_rdata_i_27_, data_rdata_i_26_, data_rdata_i_25_, data_rdata_i_24_, data_rdata_i_23_, data_rdata_i_22_, data_rdata_i_21_, data_rdata_i_20_, data_rdata_i_19_, data_rdata_i_18_, data_rdata_i_17_, data_rdata_i_16_, data_rdata_i_15_, data_rdata_i_14_, data_rdata_i_13_, data_rdata_i_12_, data_rdata_i_11_, data_rdata_i_10_, data_rdata_i_9_, data_rdata_i_8_, data_rdata_i_7_, data_rdata_i_6_, data_rdata_i_5_, data_rdata_i_4_, data_rdata_i_3_, data_rdata_i_2_, data_rdata_i_1_, data_rdata_i_0_, data_err_i, dummy_instr_id_o, rf_raddr_a_o_4_, rf_raddr_a_o_3_, rf_raddr_a_o_2_, rf_raddr_a_o_1_, rf_raddr_a_o_0_, rf_raddr_b_o_4_, rf_raddr_b_o_3_, rf_raddr_b_o_2_, rf_raddr_b_o_1_, rf_raddr_b_o_0_, rf_waddr_wb_o_4_, rf_waddr_wb_o_3_, rf_waddr_wb_o_2_, rf_waddr_wb_o_1_, rf_waddr_wb_o_0_, rf_we_wb_o, rf_wdata_wb_ecc_o_31_, rf_wdata_wb_ecc_o_30_, rf_wdata_wb_ecc_o_29_, rf_wdata_wb_ecc_o_28_, rf_wdata_wb_ecc_o_27_, rf_wdata_wb_ecc_o_26_, rf_wdata_wb_ecc_o_25_, rf_wdata_wb_ecc_o_24_, rf_wdata_wb_ecc_o_23_, rf_wdata_wb_ecc_o_22_, rf_wdata_wb_ecc_o_21_, rf_wdata_wb_ecc_o_20_, rf_wdata_wb_ecc_o_19_, rf_wdata_wb_ecc_o_18_, rf_wdata_wb_ecc_o_17_, rf_wdata_wb_ecc_o_16_, rf_wdata_wb_ecc_o_15_, rf_wdata_wb_ecc_o_14_, rf_wdata_wb_ecc_o_13_, rf_wdata_wb_ecc_o_12_, rf_wdata_wb_ecc_o_11_, rf_wdata_wb_ecc_o_10_, rf_wdata_wb_ecc_o_9_, rf_wdata_wb_ecc_o_8_, rf_wdata_wb_ecc_o_7_, rf_wdata_wb_ecc_o_6_, rf_wdata_wb_ecc_o_5_, rf_wdata_wb_ecc_o_4_, rf_wdata_wb_ecc_o_3_, rf_wdata_wb_ecc_o_2_, rf_wdata_wb_ecc_o_1_, rf_wdata_wb_ecc_o_0_, rf_rdata_a_ecc_i_31_, rf_rdata_a_ecc_i_30_, rf_rdata_a_ecc_i_29_, rf_rdata_a_ecc_i_28_, rf_rdata_a_ecc_i_27_, rf_rdata_a_ecc_i_26_, rf_rdata_a_ecc_i_25_, rf_rdata_a_ecc_i_24_, rf_rdata_a_ecc_i_23_, rf_rdata_a_ecc_i_22_, rf_rdata_a_ecc_i_21_, rf_rdata_a_ecc_i_20_, rf_rdata_a_ecc_i_19_, rf_rdata_a_ecc_i_18_, rf_rdata_a_ecc_i_17_, rf_rdata_a_ecc_i_16_, rf_rdata_a_ecc_i_15_, rf_rdata_a_ecc_i_14_, rf_rdata_a_ecc_i_13_, rf_rdata_a_ecc_i_12_, rf_rdata_a_ecc_i_11_, rf_rdata_a_ecc_i_10_, rf_rdata_a_ecc_i_9_, rf_rdata_a_ecc_i_8_, rf_rdata_a_ecc_i_7_, rf_rdata_a_ecc_i_6_, rf_rdata_a_ecc_i_5_, rf_rdata_a_ecc_i_4_, rf_rdata_a_ecc_i_3_, rf_rdata_a_ecc_i_2_, rf_rdata_a_ecc_i_1_, rf_rdata_a_ecc_i_0_, rf_rdata_b_ecc_i_31_, rf_rdata_b_ecc_i_30_, rf_rdata_b_ecc_i_29_, rf_rdata_b_ecc_i_28_, rf_rdata_b_ecc_i_27_, rf_rdata_b_ecc_i_26_, rf_rdata_b_ecc_i_25_, rf_rdata_b_ecc_i_24_, rf_rdata_b_ecc_i_23_, rf_rdata_b_ecc_i_22_, rf_rdata_b_ecc_i_21_, rf_rdata_b_ecc_i_20_, rf_rdata_b_ecc_i_19_, rf_rdata_b_ecc_i_18_, rf_rdata_b_ecc_i_17_, rf_rdata_b_ecc_i_16_, rf_rdata_b_ecc_i_15_, rf_rdata_b_ecc_i_14_, rf_rdata_b_ecc_i_13_, rf_rdata_b_ecc_i_12_, rf_rdata_b_ecc_i_11_, rf_rdata_b_ecc_i_10_, rf_rdata_b_ecc_i_9_, rf_rdata_b_ecc_i_8_, rf_rdata_b_ecc_i_7_, rf_rdata_b_ecc_i_6_, rf_rdata_b_ecc_i_5_, rf_rdata_b_ecc_i_4_, rf_rdata_b_ecc_i_3_, rf_rdata_b_ecc_i_2_, rf_rdata_b_ecc_i_1_, rf_rdata_b_ecc_i_0_, ic_tag_req_o_1_, ic_tag_req_o_0_, ic_tag_write_o, ic_tag_addr_o_7_, ic_tag_addr_o_6_, ic_tag_addr_o_5_, ic_tag_addr_o_4_, ic_tag_addr_o_3_, ic_tag_addr_o_2_, ic_tag_addr_o_1_, ic_tag_addr_o_0_, ic_tag_wdata_o_21_, ic_tag_wdata_o_20_, ic_tag_wdata_o_19_, ic_tag_wdata_o_18_, ic_tag_wdata_o_17_, ic_tag_wdata_o_16_, ic_tag_wdata_o_15_, ic_tag_wdata_o_14_, ic_tag_wdata_o_13_, ic_tag_wdata_o_12_, ic_tag_wdata_o_11_, ic_tag_wdata_o_10_, ic_tag_wdata_o_9_, ic_tag_wdata_o_8_, ic_tag_wdata_o_7_, ic_tag_wdata_o_6_, ic_tag_wdata_o_5_, ic_tag_wdata_o_4_, ic_tag_wdata_o_3_, ic_tag_wdata_o_2_, ic_tag_wdata_o_1_, ic_tag_wdata_o_0_, ic_tag_rdata_i_43_, ic_tag_rdata_i_42_, ic_tag_rdata_i_41_, ic_tag_rdata_i_40_, ic_tag_rdata_i_39_, ic_tag_rdata_i_38_, ic_tag_rdata_i_37_, ic_tag_rdata_i_36_, ic_tag_rdata_i_35_, ic_tag_rdata_i_34_, ic_tag_rdata_i_33_, ic_tag_rdata_i_32_, ic_tag_rdata_i_31_, ic_tag_rdata_i_30_, ic_tag_rdata_i_29_, ic_tag_rdata_i_28_, ic_tag_rdata_i_27_, ic_tag_rdata_i_26_, ic_tag_rdata_i_25_, ic_tag_rdata_i_24_, ic_tag_rdata_i_23_, ic_tag_rdata_i_22_, ic_tag_rdata_i_21_, ic_tag_rdata_i_20_, ic_tag_rdata_i_19_, ic_tag_rdata_i_18_, ic_tag_rdata_i_17_, ic_tag_rdata_i_16_, ic_tag_rdata_i_15_, ic_tag_rdata_i_14_, ic_tag_rdata_i_13_, ic_tag_rdata_i_12_, ic_tag_rdata_i_11_, ic_tag_rdata_i_10_, ic_tag_rdata_i_9_, ic_tag_rdata_i_8_, ic_tag_rdata_i_7_, ic_tag_rdata_i_6_, ic_tag_rdata_i_5_, ic_tag_rdata_i_4_, ic_tag_rdata_i_3_, ic_tag_rdata_i_2_, ic_tag_rdata_i_1_, ic_tag_rdata_i_0_, ic_data_req_o_1_, ic_data_req_o_0_, ic_data_write_o, ic_data_addr_o_7_, ic_data_addr_o_6_, ic_data_addr_o_5_, ic_data_addr_o_4_, ic_data_addr_o_3_, ic_data_addr_o_2_, ic_data_addr_o_1_, ic_data_addr_o_0_, ic_data_wdata_o_63_, ic_data_wdata_o_62_, ic_data_wdata_o_61_, ic_data_wdata_o_60_, ic_data_wdata_o_59_, ic_data_wdata_o_58_, ic_data_wdata_o_57_, ic_data_wdata_o_56_, ic_data_wdata_o_55_, ic_data_wdata_o_54_, ic_data_wdata_o_53_, ic_data_wdata_o_52_, ic_data_wdata_o_51_, ic_data_wdata_o_50_, ic_data_wdata_o_49_, ic_data_wdata_o_48_, ic_data_wdata_o_47_, ic_data_wdata_o_46_, ic_data_wdata_o_45_, ic_data_wdata_o_44_, ic_data_wdata_o_43_, ic_data_wdata_o_42_, ic_data_wdata_o_41_, ic_data_wdata_o_40_, ic_data_wdata_o_39_, ic_data_wdata_o_38_, ic_data_wdata_o_37_, ic_data_wdata_o_36_, ic_data_wdata_o_35_, ic_data_wdata_o_34_, ic_data_wdata_o_33_, ic_data_wdata_o_32_, ic_data_wdata_o_31_, ic_data_wdata_o_30_, ic_data_wdata_o_29_, ic_data_wdata_o_28_, ic_data_wdata_o_27_, ic_data_wdata_o_26_, ic_data_wdata_o_25_, ic_data_wdata_o_24_, ic_data_wdata_o_23_, ic_data_wdata_o_22_, ic_data_wdata_o_21_, ic_data_wdata_o_20_, ic_data_wdata_o_19_, ic_data_wdata_o_18_, ic_data_wdata_o_17_, ic_data_wdata_o_16_, ic_data_wdata_o_15_, ic_data_wdata_o_14_, ic_data_wdata_o_13_, ic_data_wdata_o_12_, ic_data_wdata_o_11_, ic_data_wdata_o_10_, ic_data_wdata_o_9_, ic_data_wdata_o_8_, ic_data_wdata_o_7_, ic_data_wdata_o_6_, ic_data_wdata_o_5_, ic_data_wdata_o_4_, ic_data_wdata_o_3_, ic_data_wdata_o_2_, ic_data_wdata_o_1_, ic_data_wdata_o_0_, ic_data_rdata_i_127_, ic_data_rdata_i_126_, ic_data_rdata_i_125_, ic_data_rdata_i_124_, ic_data_rdata_i_123_, ic_data_rdata_i_122_, ic_data_rdata_i_121_, ic_data_rdata_i_120_, ic_data_rdata_i_119_, ic_data_rdata_i_118_, ic_data_rdata_i_117_, ic_data_rdata_i_116_, ic_data_rdata_i_115_, ic_data_rdata_i_114_, ic_data_rdata_i_113_, ic_data_rdata_i_112_, ic_data_rdata_i_111_, ic_data_rdata_i_110_, ic_data_rdata_i_109_, ic_data_rdata_i_108_, ic_data_rdata_i_107_, ic_data_rdata_i_106_, ic_data_rdata_i_105_, ic_data_rdata_i_104_, ic_data_rdata_i_103_, ic_data_rdata_i_102_, ic_data_rdata_i_101_, ic_data_rdata_i_100_, ic_data_rdata_i_99_, ic_data_rdata_i_98_, ic_data_rdata_i_97_, ic_data_rdata_i_96_, ic_data_rdata_i_95_, ic_data_rdata_i_94_, ic_data_rdata_i_93_, ic_data_rdata_i_92_, ic_data_rdata_i_91_, ic_data_rdata_i_90_, ic_data_rdata_i_89_, ic_data_rdata_i_88_, ic_data_rdata_i_87_, ic_data_rdata_i_86_, ic_data_rdata_i_85_, ic_data_rdata_i_84_, ic_data_rdata_i_83_, ic_data_rdata_i_82_, ic_data_rdata_i_81_, ic_data_rdata_i_80_, ic_data_rdata_i_79_, ic_data_rdata_i_78_, ic_data_rdata_i_77_, ic_data_rdata_i_76_, ic_data_rdata_i_75_, ic_data_rdata_i_74_, ic_data_rdata_i_73_, ic_data_rdata_i_72_, ic_data_rdata_i_71_, ic_data_rdata_i_70_, ic_data_rdata_i_69_, ic_data_rdata_i_68_, ic_data_rdata_i_67_, ic_data_rdata_i_66_, ic_data_rdata_i_65_, ic_data_rdata_i_64_, ic_data_rdata_i_63_, ic_data_rdata_i_62_, ic_data_rdata_i_61_, ic_data_rdata_i_60_, ic_data_rdata_i_59_, ic_data_rdata_i_58_, ic_data_rdata_i_57_, ic_data_rdata_i_56_, ic_data_rdata_i_55_, ic_data_rdata_i_54_, ic_data_rdata_i_53_, ic_data_rdata_i_52_, ic_data_rdata_i_51_, ic_data_rdata_i_50_, ic_data_rdata_i_49_, ic_data_rdata_i_48_, ic_data_rdata_i_47_, ic_data_rdata_i_46_, ic_data_rdata_i_45_, ic_data_rdata_i_44_, ic_data_rdata_i_43_, ic_data_rdata_i_42_, ic_data_rdata_i_41_, ic_data_rdata_i_40_, ic_data_rdata_i_39_, ic_data_rdata_i_38_, ic_data_rdata_i_37_, ic_data_rdata_i_36_, ic_data_rdata_i_35_, ic_data_rdata_i_34_, ic_data_rdata_i_33_, ic_data_rdata_i_32_, ic_data_rdata_i_31_, ic_data_rdata_i_30_, ic_data_rdata_i_29_, ic_data_rdata_i_28_, ic_data_rdata_i_27_, ic_data_rdata_i_26_, ic_data_rdata_i_25_, ic_data_rdata_i_24_, ic_data_rdata_i_23_, ic_data_rdata_i_22_, ic_data_rdata_i_21_, ic_data_rdata_i_20_, ic_data_rdata_i_19_, ic_data_rdata_i_18_, ic_data_rdata_i_17_, ic_data_rdata_i_16_, ic_data_rdata_i_15_, ic_data_rdata_i_14_, ic_data_rdata_i_13_, ic_data_rdata_i_12_, ic_data_rdata_i_11_, ic_data_rdata_i_10_, ic_data_rdata_i_9_, ic_data_rdata_i_8_, ic_data_rdata_i_7_, ic_data_rdata_i_6_, ic_data_rdata_i_5_, ic_data_rdata_i_4_, ic_data_rdata_i_3_, ic_data_rdata_i_2_, ic_data_rdata_i_1_, ic_data_rdata_i_0_, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i_14_, irq_fast_i_13_, irq_fast_i_12_, irq_fast_i_11_, irq_fast_i_10_, irq_fast_i_9_, irq_fast_i_8_, irq_fast_i_7_, irq_fast_i_6_, irq_fast_i_5_, irq_fast_i_4_, irq_fast_i_3_, irq_fast_i_2_, irq_fast_i_1_, irq_fast_i_0_, irq_nm_i, irq_pending_o, debug_req_i, crash_dump_o_127_, crash_dump_o_126_, crash_dump_o_125_, crash_dump_o_124_, crash_dump_o_123_, crash_dump_o_122_, crash_dump_o_121_, crash_dump_o_120_, crash_dump_o_119_, crash_dump_o_118_, crash_dump_o_117_, crash_dump_o_116_, crash_dump_o_115_, crash_dump_o_114_, crash_dump_o_113_, crash_dump_o_112_, crash_dump_o_111_, crash_dump_o_110_, crash_dump_o_109_, crash_dump_o_108_, crash_dump_o_107_, crash_dump_o_106_, crash_dump_o_105_, crash_dump_o_104_, crash_dump_o_103_, crash_dump_o_102_, crash_dump_o_101_, crash_dump_o_100_, crash_dump_o_99_, crash_dump_o_98_, crash_dump_o_97_, crash_dump_o_96_, crash_dump_o_95_, crash_dump_o_94_, crash_dump_o_93_, crash_dump_o_92_, crash_dump_o_91_, crash_dump_o_90_, crash_dump_o_89_, crash_dump_o_88_, crash_dump_o_87_, crash_dump_o_86_, crash_dump_o_85_, crash_dump_o_84_, crash_dump_o_83_, crash_dump_o_82_, crash_dump_o_81_, crash_dump_o_80_, crash_dump_o_79_, crash_dump_o_78_, crash_dump_o_77_, crash_dump_o_76_, crash_dump_o_75_, crash_dump_o_74_, crash_dump_o_73_, crash_dump_o_72_, crash_dump_o_71_, crash_dump_o_70_, crash_dump_o_69_, crash_dump_o_68_, crash_dump_o_67_, crash_dump_o_66_, crash_dump_o_65_, crash_dump_o_64_, crash_dump_o_63_, crash_dump_o_62_, crash_dump_o_61_, crash_dump_o_60_, crash_dump_o_59_, crash_dump_o_58_, crash_dump_o_57_, crash_dump_o_56_, crash_dump_o_55_, crash_dump_o_54_, crash_dump_o_53_, crash_dump_o_52_, crash_dump_o_51_, crash_dump_o_50_, crash_dump_o_49_, crash_dump_o_48_, crash_dump_o_47_, crash_dump_o_46_, crash_dump_o_45_, crash_dump_o_44_, crash_dump_o_43_, crash_dump_o_42_, crash_dump_o_41_, crash_dump_o_40_, crash_dump_o_39_, crash_dump_o_38_, crash_dump_o_37_, crash_dump_o_36_, crash_dump_o_35_, crash_dump_o_34_, crash_dump_o_33_, crash_dump_o_32_, crash_dump_o_31_, crash_dump_o_30_, crash_dump_o_29_, crash_dump_o_28_, crash_dump_o_27_, crash_dump_o_26_, crash_dump_o_25_, crash_dump_o_24_, crash_dump_o_23_, crash_dump_o_22_, crash_dump_o_21_, crash_dump_o_20_, crash_dump_o_19_, crash_dump_o_18_, crash_dump_o_17_, crash_dump_o_16_, crash_dump_o_15_, crash_dump_o_14_, crash_dump_o_13_, crash_dump_o_12_, crash_dump_o_11_, crash_dump_o_10_, crash_dump_o_9_, crash_dump_o_8_, crash_dump_o_7_, crash_dump_o_6_, crash_dump_o_5_, crash_dump_o_4_, crash_dump_o_3_, crash_dump_o_2_, crash_dump_o_1_, crash_dump_o_0_, fetch_enable_i, alert_minor_o, alert_major_o, core_busy_o , n15981, n15965, n15980, n15964, n15985, n15963, n16056, n15962, n16055, n15961, n15984, n15960, n16054, n15959, n15983, n15958, n15990, n15957, n15989, n15956, n15988, n15955, n16053, n15954, n15987, n15953, n15986, n15952, n15995, n15951, n16052, n15950, n15994, n15949, n15993, n15948, n15992, n15947, n15991, n15946, n16051, n15945, n15996, n15944, n15999, n15943, n15998, n15942, n16002, n15941, n15997, n15940, n16007, n15939, n15936, n15938, n15935, n16126, n15934, n15937, n10609, n15933, n15978, cs_registers_i_mhpmcounter_0__63_, n10614, n10616, n10618, n10619, n10620, n10624, cs_registers_i_mhpmcounter_0__29_, cs_registers_i_mhpmcounter_0__61_, cs_registers_i_mhpmcounter_2__63_, cs_registers_i_mhpmcounter_2__62_, cs_registers_i_mhpmcounter_2__61_, n10630, n10634, cs_registers_i_mhpmcounter_0__28_, cs_registers_i_mhpmcounter_0__60_, cs_registers_i_mhpmcounter_2__28_, n10638, n10639, n10640, n10641, n10642, n10643, instr_fetch_err_plus2, n10645, n10649, cs_registers_i_mhpmcounter_0__17_, cs_registers_i_mhpmcounter_0__49_, cs_registers_i_mhpmcounter_2__17_, cs_registers_i_mhpmcounter_2__49_, n16029, n16196, n10656, n10657, n15975, n10659, n10660, n10664, cs_registers_i_mhpmcounter_0__0_, cs_registers_i_mhpmcounter_0__1_, cs_registers_i_mhpmcounter_0__2_, n10668, n10672, cs_registers_i_mhpmcounter_0__35_, cs_registers_i_mhpmcounter_2__35_, cs_registers_i_mhpmcounter_2__3_, n10676, n16050, n10678, n10682, cs_registers_i_mhpmcounter_0__39_, cs_registers_i_mhpmcounter_0__7_, cs_registers_i_mhpmcounter_2__39_, cs_registers_i_mhpmcounter_2__7_, n10687, n10688, n15974, n10690, n15932, n15977, cs_registers_i_mhpmcounter_0__36_, cs_registers_i_mhpmcounter_0__4_, cs_registers_i_mhpmcounter_2__36_, cs_registers_i_mhpmcounter_2__4_, n10697, n10699, n10700, n10701, n10702, n10703, cs_registers_i_mhpmcounter_0__38_, cs_registers_i_mhpmcounter_0__6_, cs_registers_i_mhpmcounter_2__38_, cs_registers_i_mhpmcounter_2__6_, n10710, n10712, n16005, n10714, n10715, n10716, cs_registers_i_mhpmcounter_0__40_, cs_registers_i_mhpmcounter_0__8_, cs_registers_i_mhpmcounter_2__40_, cs_registers_i_mhpmcounter_2__8_, n16023, n10724, n10726, n10727, n10728, n10729, n10730, cs_registers_i_mhpmcounter_0__41_, cs_registers_i_mhpmcounter_0__9_, cs_registers_i_mhpmcounter_2__41_, cs_registers_i_mhpmcounter_2__9_, n16039, n10738, n10740, n16022, n10742, n10743, n10744, cs_registers_i_mhpmcounter_0__10_, cs_registers_i_mhpmcounter_0__42_, cs_registers_i_mhpmcounter_2__10_, cs_registers_i_mhpmcounter_2__42_, n16024, n10752, n10754, n16021, n10756, n10757, n10758, cs_registers_i_mhpmcounter_0__11_, cs_registers_i_mhpmcounter_0__43_, cs_registers_i_mhpmcounter_2__11_, cs_registers_i_mhpmcounter_2__43_, n16133, n10767, n10771, cs_registers_i_mhpmcounter_0__12_, cs_registers_i_mhpmcounter_0__44_, cs_registers_i_mhpmcounter_2__12_, cs_registers_i_mhpmcounter_2__44_, n16025, n10777, n11303, n10778, n10779, priv_mode_id_1, n10780, n10781, cs_registers_i_mhpmcounter_0__13_, cs_registers_i_mhpmcounter_0__45_, cs_registers_i_mhpmcounter_2__13_, cs_registers_i_mhpmcounter_2__45_, n10786, n16026, n10791, n10792, n16020, n10794, n10795, n10796, cs_registers_i_mhpmcounter_0__14_, cs_registers_i_mhpmcounter_0__46_, cs_registers_i_mhpmcounter_2__14_, cs_registers_i_mhpmcounter_2__46_, n10801, n16027, n10806, n16019, n10808, n10809, n10810, cs_registers_i_mhpmcounter_0__15_, cs_registers_i_mhpmcounter_0__47_, cs_registers_i_mhpmcounter_2__15_, cs_registers_i_mhpmcounter_2__47_, n10815, n16028, n16043, n10821, n16018, n10823, n10824, n10825, cs_registers_i_mhpmcounter_0__16_, cs_registers_i_mhpmcounter_0__48_, cs_registers_i_mhpmcounter_2__16_, cs_registers_i_mhpmcounter_2__48_, n10830, n10834, n10835, n10836, n10837, n10838, n16017, n10840, cs_registers_i_mhpmcounter_0__18_, cs_registers_i_mhpmcounter_0__50_, cs_registers_i_mhpmcounter_2__18_, cs_registers_i_mhpmcounter_2__50_, n10845, n16030, n10850, n10851, n10852, n10853, n10854, n16049, n16006, n10857, cs_registers_i_mhpmcounter_0__19_, cs_registers_i_mhpmcounter_0__51_, cs_registers_i_mhpmcounter_2__19_, cs_registers_i_mhpmcounter_2__51_, n10862, n16031, n10867, n10868, n10869, n10870, n16012, n10872, cs_registers_i_mhpmcounter_0__20_, cs_registers_i_mhpmcounter_0__52_, cs_registers_i_mhpmcounter_2__20_, cs_registers_i_mhpmcounter_2__52_, n10877, n10881, n10882, n10883, n10884, n10885, n16013, n10887, cs_registers_i_mhpmcounter_0__22_, cs_registers_i_mhpmcounter_0__54_, cs_registers_i_mhpmcounter_2__22_, cs_registers_i_mhpmcounter_2__54_, n10892, n16033, n10897, n10898, n10899, n10900, n16003, n10902, cs_registers_i_mhpmcounter_0__23_, cs_registers_i_mhpmcounter_0__55_, cs_registers_i_mhpmcounter_2__23_, cs_registers_i_mhpmcounter_2__55_, n10907, n16034, n10912, n10913, n10914, n10915, n16010, n10917, cs_registers_i_mhpmcounter_0__24_, cs_registers_i_mhpmcounter_0__56_, cs_registers_i_mhpmcounter_2__24_, cs_registers_i_mhpmcounter_2__56_, n10922, n16035, n10927, n10928, n10929, n10930, n16009, n10932, cs_registers_i_mhpmcounter_0__25_, cs_registers_i_mhpmcounter_0__57_, cs_registers_i_mhpmcounter_2__25_, cs_registers_i_mhpmcounter_2__57_, n10937, n10941, n10942, n10943, n10944, n10945, n16000, n10947, cs_registers_i_mhpmcounter_0__26_, cs_registers_i_mhpmcounter_0__58_, cs_registers_i_mhpmcounter_2__26_, cs_registers_i_mhpmcounter_2__58_, n10952, n16036, n10957, n10958, n10959, n10960, n16001, n10962, cs_registers_i_mhpmcounter_0__27_, cs_registers_i_mhpmcounter_0__59_, cs_registers_i_mhpmcounter_2__27_, cs_registers_i_mhpmcounter_2__59_, n10967, n10971, n10972, n10973, n10974, n10975, n16004, n10977, n10978, n10980, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, nmi_mode, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n16081, n11304, n11487, n11481, n15798, n11018, n16032, n16037, n16038, n16040, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n15923, n15818, n16115, n11065, n16080, n16079, n16078, n16077, n16076, n16075, n16074, n16073, n16072, n16071, n16070, n16069, n16068, n16067, n16066, n16065, n16064, n16063, n16062, n16061, n16060, n16059, n16058, n16057, n10547, n10546, n15911, n15822, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n15973, n11108, n15976, n11110, n11111, n11112, n11113, cs_registers_i_mhpmcounter_0__21_, cs_registers_i_mhpmcounter_0__30_, cs_registers_i_mhpmcounter_0__32_, cs_registers_i_mhpmcounter_0__33_, cs_registers_i_mhpmcounter_0__34_, cs_registers_i_mhpmcounter_0__37_, cs_registers_i_mhpmcounter_0__53_, cs_registers_i_mhpmcounter_0__5_, cs_registers_i_mhpmcounter_2__1_, cs_registers_i_mhpmcounter_2__21_, cs_registers_i_mhpmcounter_2__2_, cs_registers_i_mhpmcounter_2__30_, cs_registers_i_mhpmcounter_2__31_, cs_registers_i_mhpmcounter_2__32_, cs_registers_i_mhpmcounter_2__33_, cs_registers_i_mhpmcounter_2__34_, cs_registers_i_mhpmcounter_2__37_, cs_registers_i_mhpmcounter_2__53_, cs_registers_i_mhpmcounter_2__5_, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n16015, n16016, n16127, n16008, n16011, n11149, n11150, n11151, n11152, n16125, n15931, n15930, n16114, n15906, n15905, n15904, n15903, n15902, n15901, n15900, n15899, n15898, n15886, n16194, n16193, n15875, n15874, n15873, n15872, n15871, n15870, n15869, n15868, n15867, n15866, n15865, n15864, n15863, n15862, n15861, n15883, n15882, n15881, n15880, n15897, n16192, n16191, n16190, n16189, n16188, n16187, n16186, n16185, n16184, n16183, n16182, n16181, n16180, n16179, n16178, n16177, n16176, n16175, n16174, n16173, n16172, n16153, n16152, n16151, n16150, n16149, n16148, n16147, n16146, n15891, n15896, n11219, n16171, n16170, n16169, n16113, n16112, n16111, n16110, n16109, n16108, n16107, n16106, n16168, n16105, n16104, n16103, n16102, n16101, n16100, n16099, n16098, n16097, n16096, n16167, n16095, n16041, n16144, n16143, n16142, n16141, n16140, n16139, n16138, ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_4, ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_3, ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_2, ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_1, ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_0, n15887, n16166, n16165, n16164, n16094, n16093, n16163, n16162, n16161, n16160, n16159, n16158, n16120, n16092, n16091, n16090, n16089, n16088, n16157, n16087, n16086, n16156, n16155, n16154, n16085, n16084, n16137, n16122, n16083, n16136, n16135, n16134, n16121, n15877, n15888, n16197, n15916, n16131, n15925, n16130, n15825, n16145, n15922, n15823, n15915, id_stage_i_controller_i_enter_debug_mode_prio_q, id_stage_i_controller_i_do_single_step_q, n15909, n15813, n15819, n16042, n15907, n10545, n10548, priv_mode_id_0, n11305, n11306, n15800, n11309, n11476, n11310, n15893, n15858, n11314, n15918, n16119, n15924, n15814, n15884, n15810, n15879, n15912, n15895, n15799, n15917, n15816, n15807, n15908, n15876, n15910, n15804, n15859, n15805, n15914, n15824, n15860, n15815, n15827, n15982, n16128, n15892, n11341, n15921, n11343, n15820, n15894, n11346, n15821, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11461, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11520, n15970, n16044, n11377, n11378, n11379, n15969, n11381, n11382, n15968, n11384, n11462, n11385, n11386, n11387, n15967, n15966, n11390, n16124, n16118, n11393, n16046, n11395, n15972, n16045, n11398, n15971, n16116, n11401, n11402, n11403, n11404, n11405, n16117, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n15812, n15803, n15793, n11463, n11468, n16132, n11470, n15929, n15878, n15920, n11472, n15927, n11477, cs_registers_i_mhpmcounter_0__3_, n15979, cs_registers_i_mhpmcounter_2__0_, n15926, n16047, n16129, n11484, n11486, n16048, n16014, cs_registers_i_mhpmcounter_2__60_, cs_registers_i_mhpmcounter_2__29_, n11494, n11497, n16195, n10765, n11507, cs_registers_i_mhpmcounter_0__62_, cs_registers_i_mhpmcounter_0__31_, n11511, n11518, n11521, n14858, n15022, n15310, n15145, n15259, n14806, n15044, n15194, n15165, n15578, n15102, n15419, n14828, n15752, n15049, n14962, n15305, n15553, n14984, n14994, n15075, n15337, n14889, n15120, n15333, n15656, n14981, n15146, n15642, n15085, n15089, n15162, n15300, n15711, n15453, n14867, n15359, n15696, n14955, n15101, n14844, n14997, n15313, n15495, n15598, n15076, n14813, n14894, n15509, n15096, n15543, n15549, n15732, n15399, n15540, n14810, n15209, n15647, n15702, n15555, n14931, n15295, n15195, n15319, n15452, n15173, n15779, n15363, n15500, n14795, n14912, n15180, n15528, n15311, n15216, n15439, n15464, n15105, n15427, n15738, n15035, n15286, n15742, n15253, n14939, n15348, n15535, n15449, n15245, n15671, n15255, n15139, n15274, n15579, n15434, n15352, n15334, n15007, n14978, n15715, n15230, n15457, n14857, n14871, n15095, n15005, n15367, n15382, n15210, n15402, n15629, n15126, n15001, n14824, n15289, n15624, n15615, n15755, n15753, n15197, n15583, n15408, n14869, n15386, n15155, n15531, n14950, n14959, n15090, n14907, n15061, n15567, n15584, n15680, n15377, n14974, n15364, n15397, n15657, n15706, n15610, n14905, n14996, n15028, n14930, n14964, n15018, n15002, n15666, n15699, n15083, n15281, n15082, n15136, n15390, n15396, n15668, n15144, n15569, n15237, n15485, n15737, n15762, n14802, n15107, n15674, n15203, n14926, n15700, n15128, n15763, n15443, n15631, n14929, n15678, n14899, n14911, n15006, n15284, n15297, n15694, n14918, n15264, n15244, n14897, n15034, n15338, n15053, n15117, n14881, n15213, n15123, n14944, n14975, n14801, n15461, n15356, n15030, n15058, n15436, n15703, n14972, n15276, n14812, n15529, n15676, n15254, n15488, n15565, n15079, n15772, n15635, n15458, n15133, n14993, n15198, n15234, n15783, n14831, n14854, n15070, n15186, n15669, n14841, n15655, n14816, n15721, n15777, n15008, n15009, n15039, n15534, n15438, n15557, n15329, n15292, n15603, n15758, n15645, n15560, n15100, n15731, n15767, n15004, n15068, n15059, n15243, n14951, n14830, n14794, n14901, n15369, n15116, n14970, n15413, n15526, n15476, n15091, n14792, n15312, n15403, n20894, n14935, n15564, n14922, n15723, n14908, n15539, n15612, n15520, n14868, n15507, n15024, n15094, n15646, n15071, n15472, n15287, n15012, n14875, n15092, n15221, n15261, n14878, n14843, n15063, n15505, n15527, n14840, n15684, n14838, n14865, n15681, n15558, n15391, n15351, n15563, n15045, n15097, n15229, n15317, n14800, n14803, n15484, n15219, n15185, n14882, n14827, n15335, n15459, n15513, n14913, n15157, n15478, n15545, n15099, n15160, n15395, n15316, n15379, n14851, n15775, n15542, n15613, n15191, n14872, n15582, n15764, n14988, n15704, n15770, n14823, n14814, n15471, n14817, n15376, n15258, n15052, n15639, n15765, n15291, n14876, n15188, n14917, n15381, n15416, n15087, n15371, n14808, n15062, n15538, n15698, n14958, n14826, n15228, n15760, n15013, n15246, n15130, n14973, n15385, n15410, n15027, n15415, n15514, n15278, n15033, n15400, n15423, n15517, n15345, n15301, n15781, n14825, n14921, n15113, n15304, n15622, n15620, n15486, n15498, n14938, n15588, n15277, n15242, n14864, n15283, n15321, n14859, n15177, n15554, n14885, n15435, n15648, n15153, n15709, n15282, n15437, n14999, n14799, n15467, n15548, n14804, n15241, n15720, n15134, n15406, n15456, n15586, n15651, n15688, n15362, n15743, n14797, n15215, n15633, n15510, n15019, n15572, n15341, n14880, n15773, n15469, n14989, n14998, n15183, n14941, n15078, n14822, n15148, n14942, n14990, n15468, n15129, n15235, n15477, n15734, n15231, n15710, n15636, n15201, n15626, n15315, n15728, n15644, n15273, n15205, n15239, n15298, n15294, n15414, n15649, n14874, n15643, n15675, n15025, n15733, n15374, n15713, n15494, n15223, n15663, n15550, n15530, n15673, n14916, n15288, n15296, n15330, n15121, n14957, n15141, n15306, n15614, n15693, n15716, n15761, n14956, n15735, n15232, n15200, n15060, n15571, n14960, n15621, n15072, n15174, n15451, n15159, n14818, n15618, n14948, n14850, n15346, n14952, n15503, n15279, n15178, n14967, n15522, n15263, n15533, n14963, n14842, n15041, n15577, n14992, n15506, n14853, n15780, n14852, n15236, n15532, n15428, n15179, n15418, n15450, n15115, n14979, n15591, n15354, n14886, n14892, n15623, n15559, n14968, n15320, n15175, n15525, n15653, n15110, n15192, n14919, n14821, n15574, n14947, n15048, n15014, n15168, n15344, n14811, n15054, n15166, n15260, n15608, n15508, n15405, n14820, n14928, n15566, n14903, n14891, n15616, n15147, n15524, n14927, n15073, n14923, n15328, n15609, n15705, n15782, n14914, n15055, n15754, n14896, n15679, n15164, n15086, n15501, n14848, n15124, n15685, n15491, n15015, n15140, n15360, n15474, n15740, n14796, n15190, n15447, n15098, n14870, n14977, n15302, n15023, n14982, n15046, n15339, n15718, n15430, n14835, n15189, n15251, n15778, n15383, n15003, n15431, n15512, n15275, n15463, n15421, n15519, n15161, n15355, n15561, n15208, n14863, n15714, n15749, n15759, n15632, n15365, n15747, n14860, n15156, n15187, n15604, n15336, n15375, n15342, n15404, n15257, n15118, n15499, n15585, n15575, n15619, n15163, n15701, n15465, n15167, n15268, n15370, n15487, n15220, n15088, n15309, n15521, n15625, n14845, n14856, n14887, n15067, n15470, n15768, n15171, n15446, n15248, n15687, n15412, n15043, n15104, n14890, n14936, n15247, n14991, n15384, n15690, n14834, n15717, n14966, n15448, n15432, n15659, n15686, n15212, n15020, n15303, n15214, n15314, n15181, n15047, n15154, n15401, n14862, n14980, n15318, n15589, n14924, n15462, n15016, n14940, n15358, n15409, n14829, n14920, n15712, n15460, n14866, n15143, n14832, n14855, n15466, n14847, n15056, n15637, n15660, n15597, n15125, n14805, n15069, n15581, n15724, n15211, n15222, n15066, n15176, n15592, n15158, n15373, n15601, n15748, n14888, n15587, n15349, n15350, n14949, n14971, n15372, n15599, n14983, n15347, n15380, n15650, n15727, n14877, n15325, n15324, n15119, n15106, n15407, n15233, n15691, n14833, n15745, n15327, n14986, n15425, n15149, n15602, n15692, n15658, n15207, n14807, n15594, n15766, n14879, n15111, n15475, n15152, n15299, n14965, n15455, n15667, n15093, n15326, n15249, n15074, n15661, n15473, n15172, n15388, n15000, n15227, n15114, n15366, n15307, n15689, n14861, n15638, n15184, n15593, n14809, n15280, n15017, n14849, n15193, n14987, n15265, n14898, n14925, n15109, n15011, n15270, n15562, n15739, n15196, n15708, n14895, n15741, n15677, n15670, n15672, n15323, n15511, n15695, n15361, n15537, n15634, n15081, n15202, n15256, n15750, n15084, n15343, n15262, n15454, n15568, n14904, n15142, n14946, n15627, n15040, n15744, n15445, n14793, n15151, n15077, n15132, n15544, n15665, n14883, n15080, n15226, n15492, n14839, n15523, n15417, n15387, n15206, n15641, n14976, n15150, n15607, n15751, n15340, n14954, n15444, n15021, n15285, n15757, n15774, n15331, n15037, n15240, n15730, n15489, n15722, n15606, n15010, n15424, n15547, n15392, n15064, n15138, n14884, n15199, n15411, n15652, n15576, n15429, n14943, n15029, n14934, n15269, n15422, n14969, n14900, n15218, n15332, n14798, n15137, n15042, n14995, n15420, n15122, n15182, n15490, n14873, n15169, n14915, n15515, n15611, n15725, n14910, n15031, n15026, n15573, n15493, n15496, n15719, n14893, n15112, n15252, n15426, n15127, n15536, n15441, n15541, n15204, n15442, n15271, n14906, n15483, n15580, n14937, n15596, n15225, n15726, n15038, n15065, n15697, n15481, n15497, n15518, n15736, n15272, n14815, n14902, n15398, n15322, n15353, n15546, n15502, n14945, n15504, n15050, n15654, n15769, n15357, n15482, n15368, n14846, n15433, n15378, n14836, n15057, n15682, n14909, n15516, n15266, n15628, n15393, n15308, n15590, n15103, n14933, n15394, n20877, n15479, n15480, n15108, n15217, n15776, n15707, n15662, n15051, n15224, n15756, n14932, n14985, n15600, n15595, n15250, n15389, n15640, n14953, n15729, n15551, n15440, n15552, n14961, n15238, n15605, n15135, n15630, n15664, n15570, n15746, n14819, n15267, n15290, n15683, n14837, n15032, n15170, n15771, n15036, n15131, n15293, n15617);
input rst_ni, hart_id_i_31_, hart_id_i_30_, hart_id_i_29_, hart_id_i_28_, hart_id_i_27_, hart_id_i_26_, hart_id_i_25_, hart_id_i_24_, hart_id_i_23_, hart_id_i_22_, hart_id_i_21_, hart_id_i_20_, hart_id_i_19_, hart_id_i_18_, hart_id_i_17_, hart_id_i_16_, hart_id_i_15_, hart_id_i_14_, hart_id_i_13_, hart_id_i_12_, hart_id_i_11_, hart_id_i_10_, hart_id_i_9_, hart_id_i_8_, hart_id_i_7_, hart_id_i_6_, hart_id_i_5_, hart_id_i_4_, hart_id_i_3_, hart_id_i_2_, hart_id_i_1_, hart_id_i_0_, boot_addr_i_31_, boot_addr_i_30_, boot_addr_i_29_, boot_addr_i_28_, boot_addr_i_27_, boot_addr_i_26_, boot_addr_i_25_, boot_addr_i_24_, boot_addr_i_23_, boot_addr_i_22_, boot_addr_i_21_, boot_addr_i_20_, boot_addr_i_19_, boot_addr_i_18_, boot_addr_i_17_, boot_addr_i_16_, boot_addr_i_15_, boot_addr_i_14_, boot_addr_i_13_, boot_addr_i_12_, boot_addr_i_11_, boot_addr_i_10_, boot_addr_i_9_, boot_addr_i_8_, boot_addr_i_7_, boot_addr_i_6_, boot_addr_i_5_, boot_addr_i_4_, boot_addr_i_3_, boot_addr_i_2_, boot_addr_i_1_, boot_addr_i_0_, instr_gnt_i, instr_rvalid_i, instr_rdata_i_31_, instr_rdata_i_30_, instr_rdata_i_29_, instr_rdata_i_28_, instr_rdata_i_27_, instr_rdata_i_26_, instr_rdata_i_25_, instr_rdata_i_24_, instr_rdata_i_23_, instr_rdata_i_22_, instr_rdata_i_21_, instr_rdata_i_20_, instr_rdata_i_19_, instr_rdata_i_18_, instr_rdata_i_17_, instr_rdata_i_16_, instr_rdata_i_15_, instr_rdata_i_14_, instr_rdata_i_13_, instr_rdata_i_12_, instr_rdata_i_11_, instr_rdata_i_10_, instr_rdata_i_9_, instr_rdata_i_8_, instr_rdata_i_7_, instr_rdata_i_6_, instr_rdata_i_5_, instr_rdata_i_4_, instr_rdata_i_3_, instr_rdata_i_2_, instr_rdata_i_1_, instr_rdata_i_0_, instr_err_i, data_gnt_i, data_rvalid_i, data_rdata_i_31_, data_rdata_i_30_, data_rdata_i_29_, data_rdata_i_28_, data_rdata_i_27_, data_rdata_i_26_, data_rdata_i_25_, data_rdata_i_24_, data_rdata_i_23_, data_rdata_i_22_, data_rdata_i_21_, data_rdata_i_20_, data_rdata_i_19_, data_rdata_i_18_, data_rdata_i_17_, data_rdata_i_16_, data_rdata_i_15_, data_rdata_i_14_, data_rdata_i_13_, data_rdata_i_12_, data_rdata_i_11_, data_rdata_i_10_, data_rdata_i_9_, data_rdata_i_8_, data_rdata_i_7_, data_rdata_i_6_, data_rdata_i_5_, data_rdata_i_4_, data_rdata_i_3_, data_rdata_i_2_, data_rdata_i_1_, data_rdata_i_0_, data_err_i, rf_rdata_a_ecc_i_31_, rf_rdata_a_ecc_i_30_, rf_rdata_a_ecc_i_29_, rf_rdata_a_ecc_i_28_, rf_rdata_a_ecc_i_27_, rf_rdata_a_ecc_i_26_, rf_rdata_a_ecc_i_25_, rf_rdata_a_ecc_i_24_, rf_rdata_a_ecc_i_23_, rf_rdata_a_ecc_i_22_, rf_rdata_a_ecc_i_21_, rf_rdata_a_ecc_i_20_, rf_rdata_a_ecc_i_19_, rf_rdata_a_ecc_i_18_, rf_rdata_a_ecc_i_17_, rf_rdata_a_ecc_i_16_, rf_rdata_a_ecc_i_15_, rf_rdata_a_ecc_i_14_, rf_rdata_a_ecc_i_13_, rf_rdata_a_ecc_i_12_, rf_rdata_a_ecc_i_11_, rf_rdata_a_ecc_i_10_, rf_rdata_a_ecc_i_9_, rf_rdata_a_ecc_i_8_, rf_rdata_a_ecc_i_7_, rf_rdata_a_ecc_i_6_, rf_rdata_a_ecc_i_5_, rf_rdata_a_ecc_i_4_, rf_rdata_a_ecc_i_3_, rf_rdata_a_ecc_i_2_, rf_rdata_a_ecc_i_1_, rf_rdata_a_ecc_i_0_, rf_rdata_b_ecc_i_31_, rf_rdata_b_ecc_i_30_, rf_rdata_b_ecc_i_29_, rf_rdata_b_ecc_i_28_, rf_rdata_b_ecc_i_27_, rf_rdata_b_ecc_i_26_, rf_rdata_b_ecc_i_25_, rf_rdata_b_ecc_i_24_, rf_rdata_b_ecc_i_23_, rf_rdata_b_ecc_i_22_, rf_rdata_b_ecc_i_21_, rf_rdata_b_ecc_i_20_, rf_rdata_b_ecc_i_19_, rf_rdata_b_ecc_i_18_, rf_rdata_b_ecc_i_17_, rf_rdata_b_ecc_i_16_, rf_rdata_b_ecc_i_15_, rf_rdata_b_ecc_i_14_, rf_rdata_b_ecc_i_13_, rf_rdata_b_ecc_i_12_, rf_rdata_b_ecc_i_11_, rf_rdata_b_ecc_i_10_, rf_rdata_b_ecc_i_9_, rf_rdata_b_ecc_i_8_, rf_rdata_b_ecc_i_7_, rf_rdata_b_ecc_i_6_, rf_rdata_b_ecc_i_5_, rf_rdata_b_ecc_i_4_, rf_rdata_b_ecc_i_3_, rf_rdata_b_ecc_i_2_, rf_rdata_b_ecc_i_1_, rf_rdata_b_ecc_i_0_, ic_tag_rdata_i_43_, ic_tag_rdata_i_42_, ic_tag_rdata_i_41_, ic_tag_rdata_i_40_, ic_tag_rdata_i_39_, ic_tag_rdata_i_38_, ic_tag_rdata_i_37_, ic_tag_rdata_i_36_, ic_tag_rdata_i_35_, ic_tag_rdata_i_34_, ic_tag_rdata_i_33_, ic_tag_rdata_i_32_, ic_tag_rdata_i_31_, ic_tag_rdata_i_30_, ic_tag_rdata_i_29_, ic_tag_rdata_i_28_, ic_tag_rdata_i_27_, ic_tag_rdata_i_26_, ic_tag_rdata_i_25_, ic_tag_rdata_i_24_, ic_tag_rdata_i_23_, ic_tag_rdata_i_22_, ic_tag_rdata_i_21_, ic_tag_rdata_i_20_, ic_tag_rdata_i_19_, ic_tag_rdata_i_18_, ic_tag_rdata_i_17_, ic_tag_rdata_i_16_, ic_tag_rdata_i_15_, ic_tag_rdata_i_14_, ic_tag_rdata_i_13_, ic_tag_rdata_i_12_, ic_tag_rdata_i_11_, ic_tag_rdata_i_10_, ic_tag_rdata_i_9_, ic_tag_rdata_i_8_, ic_tag_rdata_i_7_, ic_tag_rdata_i_6_, ic_tag_rdata_i_5_, ic_tag_rdata_i_4_, ic_tag_rdata_i_3_, ic_tag_rdata_i_2_, ic_tag_rdata_i_1_, ic_tag_rdata_i_0_, ic_data_rdata_i_127_, ic_data_rdata_i_126_, ic_data_rdata_i_125_, ic_data_rdata_i_124_, ic_data_rdata_i_123_, ic_data_rdata_i_122_, ic_data_rdata_i_121_, ic_data_rdata_i_120_, ic_data_rdata_i_119_, ic_data_rdata_i_118_, ic_data_rdata_i_117_, ic_data_rdata_i_116_, ic_data_rdata_i_115_, ic_data_rdata_i_114_, ic_data_rdata_i_113_, ic_data_rdata_i_112_, ic_data_rdata_i_111_, ic_data_rdata_i_110_, ic_data_rdata_i_109_, ic_data_rdata_i_108_, ic_data_rdata_i_107_, ic_data_rdata_i_106_, ic_data_rdata_i_105_, ic_data_rdata_i_104_, ic_data_rdata_i_103_, ic_data_rdata_i_102_, ic_data_rdata_i_101_, ic_data_rdata_i_100_, ic_data_rdata_i_99_, ic_data_rdata_i_98_, ic_data_rdata_i_97_, ic_data_rdata_i_96_, ic_data_rdata_i_95_, ic_data_rdata_i_94_, ic_data_rdata_i_93_, ic_data_rdata_i_92_, ic_data_rdata_i_91_, ic_data_rdata_i_90_, ic_data_rdata_i_89_, ic_data_rdata_i_88_, ic_data_rdata_i_87_, ic_data_rdata_i_86_, ic_data_rdata_i_85_, ic_data_rdata_i_84_, ic_data_rdata_i_83_, ic_data_rdata_i_82_, ic_data_rdata_i_81_, ic_data_rdata_i_80_, ic_data_rdata_i_79_, ic_data_rdata_i_78_, ic_data_rdata_i_77_, ic_data_rdata_i_76_, ic_data_rdata_i_75_, ic_data_rdata_i_74_, ic_data_rdata_i_73_, ic_data_rdata_i_72_, ic_data_rdata_i_71_, ic_data_rdata_i_70_, ic_data_rdata_i_69_, ic_data_rdata_i_68_, ic_data_rdata_i_67_, ic_data_rdata_i_66_, ic_data_rdata_i_65_, ic_data_rdata_i_64_, ic_data_rdata_i_63_, ic_data_rdata_i_62_, ic_data_rdata_i_61_, ic_data_rdata_i_60_, ic_data_rdata_i_59_, ic_data_rdata_i_58_, ic_data_rdata_i_57_, ic_data_rdata_i_56_, ic_data_rdata_i_55_, ic_data_rdata_i_54_, ic_data_rdata_i_53_, ic_data_rdata_i_52_, ic_data_rdata_i_51_, ic_data_rdata_i_50_, ic_data_rdata_i_49_, ic_data_rdata_i_48_, ic_data_rdata_i_47_, ic_data_rdata_i_46_, ic_data_rdata_i_45_, ic_data_rdata_i_44_, ic_data_rdata_i_43_, ic_data_rdata_i_42_, ic_data_rdata_i_41_, ic_data_rdata_i_40_, ic_data_rdata_i_39_, ic_data_rdata_i_38_, ic_data_rdata_i_37_, ic_data_rdata_i_36_, ic_data_rdata_i_35_, ic_data_rdata_i_34_, ic_data_rdata_i_33_, ic_data_rdata_i_32_, ic_data_rdata_i_31_, ic_data_rdata_i_30_, ic_data_rdata_i_29_, ic_data_rdata_i_28_, ic_data_rdata_i_27_, ic_data_rdata_i_26_, ic_data_rdata_i_25_, ic_data_rdata_i_24_, ic_data_rdata_i_23_, ic_data_rdata_i_22_, ic_data_rdata_i_21_, ic_data_rdata_i_20_, ic_data_rdata_i_19_, ic_data_rdata_i_18_, ic_data_rdata_i_17_, ic_data_rdata_i_16_, ic_data_rdata_i_15_, ic_data_rdata_i_14_, ic_data_rdata_i_13_, ic_data_rdata_i_12_, ic_data_rdata_i_11_, ic_data_rdata_i_10_, ic_data_rdata_i_9_, ic_data_rdata_i_8_, ic_data_rdata_i_7_, ic_data_rdata_i_6_, ic_data_rdata_i_5_, ic_data_rdata_i_4_, ic_data_rdata_i_3_, ic_data_rdata_i_2_, ic_data_rdata_i_1_, ic_data_rdata_i_0_, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i_14_, irq_fast_i_13_, irq_fast_i_12_, irq_fast_i_11_, irq_fast_i_10_, irq_fast_i_9_, irq_fast_i_8_, irq_fast_i_7_, irq_fast_i_6_, irq_fast_i_5_, irq_fast_i_4_, irq_fast_i_3_, irq_fast_i_2_, irq_fast_i_1_, irq_fast_i_0_, irq_nm_i, debug_req_i, fetch_enable_i, crash_dump_o_5_, crash_dump_o_30_, crash_dump_o_21_, crash_dump_o_29_, crash_dump_o_125_, crash_dump_o_93_, crash_dump_o_28_, crash_dump_o_124_, crash_dump_o_92_, crash_dump_o_1_, crash_dump_o_17_, crash_dump_o_113_, crash_dump_o_81_, crash_dump_o_2_, crash_dump_o_98_, crash_dump_o_66_, crash_dump_o_3_, crash_dump_o_99_, crash_dump_o_67_, crash_dump_o_7_, crash_dump_o_103_, crash_dump_o_71_, crash_dump_o_4_, crash_dump_o_100_, crash_dump_o_68_, crash_dump_o_6_, crash_dump_o_102_, crash_dump_o_70_, crash_dump_o_8_, crash_dump_o_104_, crash_dump_o_72_, crash_dump_o_9_, crash_dump_o_105_, crash_dump_o_73_, crash_dump_o_10_, crash_dump_o_106_, crash_dump_o_74_, crash_dump_o_12_, crash_dump_o_108_, crash_dump_o_76_, crash_dump_o_13_, crash_dump_o_109_, crash_dump_o_77_, crash_dump_o_14_, crash_dump_o_110_, crash_dump_o_78_, crash_dump_o_15_, crash_dump_o_111_, crash_dump_o_79_, crash_dump_o_16_, crash_dump_o_112_, crash_dump_o_80_, crash_dump_o_18_, crash_dump_o_114_, crash_dump_o_82_, crash_dump_o_19_, crash_dump_o_115_, crash_dump_o_83_, crash_dump_o_20_, crash_dump_o_116_, crash_dump_o_84_, crash_dump_o_22_, crash_dump_o_118_, crash_dump_o_86_, crash_dump_o_23_, crash_dump_o_119_, crash_dump_o_87_, crash_dump_o_24_, crash_dump_o_120_, crash_dump_o_88_, crash_dump_o_25_, crash_dump_o_121_, crash_dump_o_89_, crash_dump_o_26_, crash_dump_o_122_, crash_dump_o_90_, crash_dump_o_27_, crash_dump_o_123_, crash_dump_o_91_, crash_dump_o_11_, crash_dump_o_31_, crash_dump_o_0_, crash_dump_o_33_, crash_dump_o_34_, crash_dump_o_35_, crash_dump_o_36_, crash_dump_o_37_, crash_dump_o_38_, crash_dump_o_39_, crash_dump_o_40_, crash_dump_o_41_, crash_dump_o_42_, crash_dump_o_43_, crash_dump_o_44_, crash_dump_o_45_, crash_dump_o_46_, crash_dump_o_47_, crash_dump_o_48_, crash_dump_o_49_, crash_dump_o_50_, crash_dump_o_51_, crash_dump_o_52_, crash_dump_o_53_, crash_dump_o_54_, crash_dump_o_55_, crash_dump_o_56_, crash_dump_o_57_, crash_dump_o_58_, crash_dump_o_59_, crash_dump_o_60_, crash_dump_o_61_, crash_dump_o_62_, crash_dump_o_63_, crash_dump_o_32_, crash_dump_o_107_, crash_dump_o_75_, rf_waddr_wb_o_3_, rf_waddr_wb_o_4_, rf_waddr_wb_o_2_, rf_raddr_b_o_4_, rf_raddr_a_o_4_, rf_raddr_a_o_0_, rf_raddr_a_o_2_, rf_raddr_b_o_2_, rf_raddr_a_o_1_, rf_raddr_a_o_3_, rf_raddr_b_o_0_, rf_raddr_b_o_1_, rf_raddr_b_o_3_, rf_waddr_wb_o_0_, rf_waddr_wb_o_1_, crash_dump_o_96_, crash_dump_o_97_, crash_dump_o_101_, crash_dump_o_127_, crash_dump_o_65_, crash_dump_o_117_, crash_dump_o_85_, crash_dump_o_126_, crash_dump_o_94_, crash_dump_o_95_, crash_dump_o_69_, n15981, n15965, n15980, n15964, n15985, n15963, n16056, n15962, n16055, n15961, n15984, n15960, n16054, n15959, n15983, n15958, n15990, n15957, n15989, n15956, n15988, n15955, n16053, n15954, n15987, n15953, n15986, n15952, n15995, n15951, n16052, n15950, n15994, n15949, n15993, n15948, n15992, n15947, n15991, n15946, n16051, n15945, n15996, n15944, n15999, n15943, n15998, n15942, n16002, n15941, n15997, n15940, n16007, n15939, n15936, n15938, n15935, n16126, n15934, n15937, n10609, n15933, n15978, cs_registers_i_mhpmcounter_0__63_, n10614, n10616, n10618, n10619, n10620, n10624, cs_registers_i_mhpmcounter_0__29_, cs_registers_i_mhpmcounter_0__61_, cs_registers_i_mhpmcounter_2__63_, cs_registers_i_mhpmcounter_2__62_, cs_registers_i_mhpmcounter_2__61_, n10630, n10634, cs_registers_i_mhpmcounter_0__28_, cs_registers_i_mhpmcounter_0__60_, cs_registers_i_mhpmcounter_2__28_, n10638, n10639, n10640, n10641, n10642, n10643, instr_fetch_err_plus2, n10645, n10649, cs_registers_i_mhpmcounter_0__17_, cs_registers_i_mhpmcounter_0__49_, cs_registers_i_mhpmcounter_2__17_, cs_registers_i_mhpmcounter_2__49_, n16029, n16196, n10656, n10657, n15975, n10659, n10660, n10664, cs_registers_i_mhpmcounter_0__0_, cs_registers_i_mhpmcounter_0__1_, cs_registers_i_mhpmcounter_0__2_, n10668, n10672, cs_registers_i_mhpmcounter_0__35_, cs_registers_i_mhpmcounter_2__35_, cs_registers_i_mhpmcounter_2__3_, n10676, n16050, n10678, n10682, cs_registers_i_mhpmcounter_0__39_, cs_registers_i_mhpmcounter_0__7_, cs_registers_i_mhpmcounter_2__39_, cs_registers_i_mhpmcounter_2__7_, n10687, n10688, n15974, n10690, n15932, n15977, cs_registers_i_mhpmcounter_0__36_, cs_registers_i_mhpmcounter_0__4_, cs_registers_i_mhpmcounter_2__36_, cs_registers_i_mhpmcounter_2__4_, n10697, n10699, n10700, n10701, n10702, n10703, cs_registers_i_mhpmcounter_0__38_, cs_registers_i_mhpmcounter_0__6_, cs_registers_i_mhpmcounter_2__38_, cs_registers_i_mhpmcounter_2__6_, n10710, n10712, n16005, n10714, n10715, n10716, cs_registers_i_mhpmcounter_0__40_, cs_registers_i_mhpmcounter_0__8_, cs_registers_i_mhpmcounter_2__40_, cs_registers_i_mhpmcounter_2__8_, n16023, n10724, n10726, n10727, n10728, n10729, n10730, cs_registers_i_mhpmcounter_0__41_, cs_registers_i_mhpmcounter_0__9_, cs_registers_i_mhpmcounter_2__41_, cs_registers_i_mhpmcounter_2__9_, n16039, n10738, n10740, n16022, n10742, n10743, n10744, cs_registers_i_mhpmcounter_0__10_, cs_registers_i_mhpmcounter_0__42_, cs_registers_i_mhpmcounter_2__10_, cs_registers_i_mhpmcounter_2__42_, n16024, n10752, n10754, n16021, n10756, n10757, n10758, cs_registers_i_mhpmcounter_0__11_, cs_registers_i_mhpmcounter_0__43_, cs_registers_i_mhpmcounter_2__11_, cs_registers_i_mhpmcounter_2__43_, n16133, n10767, n10771, cs_registers_i_mhpmcounter_0__12_, cs_registers_i_mhpmcounter_0__44_, cs_registers_i_mhpmcounter_2__12_, cs_registers_i_mhpmcounter_2__44_, n16025, n10777, n11303, n10778, n10779, priv_mode_id_1, n10780, n10781, cs_registers_i_mhpmcounter_0__13_, cs_registers_i_mhpmcounter_0__45_, cs_registers_i_mhpmcounter_2__13_, cs_registers_i_mhpmcounter_2__45_, n10786, n16026, n10791, n10792, n16020, n10794, n10795, n10796, cs_registers_i_mhpmcounter_0__14_, cs_registers_i_mhpmcounter_0__46_, cs_registers_i_mhpmcounter_2__14_, cs_registers_i_mhpmcounter_2__46_, n10801, n16027, n10806, n16019, n10808, n10809, n10810, cs_registers_i_mhpmcounter_0__15_, cs_registers_i_mhpmcounter_0__47_, cs_registers_i_mhpmcounter_2__15_, cs_registers_i_mhpmcounter_2__47_, n10815, n16028, n16043, n10821, n16018, n10823, n10824, n10825, cs_registers_i_mhpmcounter_0__16_, cs_registers_i_mhpmcounter_0__48_, cs_registers_i_mhpmcounter_2__16_, cs_registers_i_mhpmcounter_2__48_, n10830, n10834, n10835, n10836, n10837, n10838, n16017, n10840, cs_registers_i_mhpmcounter_0__18_, cs_registers_i_mhpmcounter_0__50_, cs_registers_i_mhpmcounter_2__18_, cs_registers_i_mhpmcounter_2__50_, n10845, n16030, n10850, n10851, n10852, n10853, n10854, n16049, n16006, n10857, cs_registers_i_mhpmcounter_0__19_, cs_registers_i_mhpmcounter_0__51_, cs_registers_i_mhpmcounter_2__19_, cs_registers_i_mhpmcounter_2__51_, n10862, n16031, n10867, n10868, n10869, n10870, n16012, n10872, cs_registers_i_mhpmcounter_0__20_, cs_registers_i_mhpmcounter_0__52_, cs_registers_i_mhpmcounter_2__20_, cs_registers_i_mhpmcounter_2__52_, n10877, n10881, n10882, n10883, n10884, n10885, n16013, n10887, cs_registers_i_mhpmcounter_0__22_, cs_registers_i_mhpmcounter_0__54_, cs_registers_i_mhpmcounter_2__22_, cs_registers_i_mhpmcounter_2__54_, n10892, n16033, n10897, n10898, n10899, n10900, n16003, n10902, cs_registers_i_mhpmcounter_0__23_, cs_registers_i_mhpmcounter_0__55_, cs_registers_i_mhpmcounter_2__23_, cs_registers_i_mhpmcounter_2__55_, n10907, n16034, n10912, n10913, n10914, n10915, n16010, n10917, cs_registers_i_mhpmcounter_0__24_, cs_registers_i_mhpmcounter_0__56_, cs_registers_i_mhpmcounter_2__24_, cs_registers_i_mhpmcounter_2__56_, n10922, n16035, n10927, n10928, n10929, n10930, n16009, n10932, cs_registers_i_mhpmcounter_0__25_, cs_registers_i_mhpmcounter_0__57_, cs_registers_i_mhpmcounter_2__25_, cs_registers_i_mhpmcounter_2__57_, n10937, n10941, n10942, n10943, n10944, n10945, n16000, n10947, cs_registers_i_mhpmcounter_0__26_, cs_registers_i_mhpmcounter_0__58_, cs_registers_i_mhpmcounter_2__26_, cs_registers_i_mhpmcounter_2__58_, n10952, n16036, n10957, n10958, n10959, n10960, n16001, n10962, cs_registers_i_mhpmcounter_0__27_, cs_registers_i_mhpmcounter_0__59_, cs_registers_i_mhpmcounter_2__27_, cs_registers_i_mhpmcounter_2__59_, n10967, n10971, n10972, n10973, n10974, n10975, n16004, n10977, n10978, n10980, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, nmi_mode, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n16081, n11304, n11487, n11481, n15798, n11018, n16032, n16037, n16038, n16040, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n15923, n15818, n16115, n11065, n16080, n16079, n16078, n16077, n16076, n16075, n16074, n16073, n16072, n16071, n16070, n16069, n16068, n16067, n16066, n16065, n16064, n16063, n16062, n16061, n16060, n16059, n16058, n16057, n10547, n10546, n15911, n15822, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n15973, n11108, n15976, n11110, n11111, n11112, n11113, cs_registers_i_mhpmcounter_0__21_, cs_registers_i_mhpmcounter_0__30_, cs_registers_i_mhpmcounter_0__32_, cs_registers_i_mhpmcounter_0__33_, cs_registers_i_mhpmcounter_0__34_, cs_registers_i_mhpmcounter_0__37_, cs_registers_i_mhpmcounter_0__53_, cs_registers_i_mhpmcounter_0__5_, cs_registers_i_mhpmcounter_2__1_, cs_registers_i_mhpmcounter_2__21_, cs_registers_i_mhpmcounter_2__2_, cs_registers_i_mhpmcounter_2__30_, cs_registers_i_mhpmcounter_2__31_, cs_registers_i_mhpmcounter_2__32_, cs_registers_i_mhpmcounter_2__33_, cs_registers_i_mhpmcounter_2__34_, cs_registers_i_mhpmcounter_2__37_, cs_registers_i_mhpmcounter_2__53_, cs_registers_i_mhpmcounter_2__5_, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n16015, n16016, n16127, n16008, n16011, n11149, n11150, n11151, n11152, n16125, n15931, n15930, n16114, n15906, n15905, n15904, n15903, n15902, n15901, n15900, n15899, n15898, n15886, n16194, n16193, n15875, n15874, n15873, n15872, n15871, n15870, n15869, n15868, n15867, n15866, n15865, n15864, n15863, n15862, n15861, n15883, n15882, n15881, n15880, n15897, n16192, n16191, n16190, n16189, n16188, n16187, n16186, n16185, n16184, n16183, n16182, n16181, n16180, n16179, n16178, n16177, n16176, n16175, n16174, n16173, n16172, n16153, n16152, n16151, n16150, n16149, n16148, n16147, n16146, n15891, n15896, n11219, n16171, n16170, n16169, n16113, n16112, n16111, n16110, n16109, n16108, n16107, n16106, n16168, n16105, n16104, n16103, n16102, n16101, n16100, n16099, n16098, n16097, n16096, n16167, n16095, n16041, n16144, n16143, n16142, n16141, n16140, n16139, n16138, ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_4, ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_3, ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_2, ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_1, ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_0, n15887, n16166, n16165, n16164, n16094, n16093, n16163, n16162, n16161, n16160, n16159, n16158, n16120, n16092, n16091, n16090, n16089, n16088, n16157, n16087, n16086, n16156, n16155, n16154, n16085, n16084, n16137, n16122, n16083, n16136, n16135, n16134, n16121, n15877, n15888, n16197, n15916, n16131, n15925, n16130, n15825, n16145, n15922, n15823, n15915, id_stage_i_controller_i_enter_debug_mode_prio_q, id_stage_i_controller_i_do_single_step_q, n15909, n15813, n15819, n16042, n15907, n10545, n10548, priv_mode_id_0, n11305, n11306, n15800, n11309, n11476, n11310, n15893, n15858, n11314, n15918, n16119, n15924, n15814, n15884, n15810, n15879, n15912, n15895, n15799, n15917, n15816, n15807, n15908, n15876, n15910, n15804, n15859, n15805, n15914, n15824, n15860, n15815, n15827, n15982, n16128, n15892, n11341, n15921, n11343, n15820, n15894, n11346, n15821, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11461, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11520, n15970, n16044, n11377, n11378, n11379, n15969, n11381, n11382, n15968, n11384, n11462, n11385, n11386, n11387, n15967, n15966, n11390, n16124, n16118, n11393, n16046, n11395, n15972, n16045, n11398, n15971, n16116, n11401, n11402, n11403, n11404, n11405, n16117, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n15812, n15803, n15793, n11463, n11468, n16132, n11470, n15929, n15878, n15920, n11472, n15927, n11477, cs_registers_i_mhpmcounter_0__3_, n15979, cs_registers_i_mhpmcounter_2__0_, n15926, n16047, n16129, n11484, n11486, n16048, n16014, cs_registers_i_mhpmcounter_2__60_, cs_registers_i_mhpmcounter_2__29_, n11494, n11497, n16195, n10765, n11507, cs_registers_i_mhpmcounter_0__62_, cs_registers_i_mhpmcounter_0__31_, n11511, n11518, n11521;
output instr_req_o, instr_addr_o_31_, instr_addr_o_30_, instr_addr_o_29_, instr_addr_o_28_, instr_addr_o_27_, instr_addr_o_26_, instr_addr_o_25_, instr_addr_o_24_, instr_addr_o_23_, instr_addr_o_22_, instr_addr_o_21_, instr_addr_o_20_, instr_addr_o_19_, instr_addr_o_18_, instr_addr_o_17_, instr_addr_o_16_, instr_addr_o_15_, instr_addr_o_14_, instr_addr_o_13_, instr_addr_o_12_, instr_addr_o_11_, instr_addr_o_10_, instr_addr_o_9_, instr_addr_o_8_, instr_addr_o_7_, instr_addr_o_6_, instr_addr_o_5_, instr_addr_o_4_, instr_addr_o_3_, instr_addr_o_2_, data_req_o, data_we_o, data_be_o_3_, data_be_o_2_, data_be_o_1_, data_be_o_0_, data_addr_o_31_, data_addr_o_30_, data_addr_o_29_, data_addr_o_28_, data_addr_o_27_, data_addr_o_26_, data_addr_o_25_, data_addr_o_24_, data_addr_o_23_, data_addr_o_22_, data_addr_o_21_, data_addr_o_20_, data_addr_o_19_, data_addr_o_18_, data_addr_o_17_, data_addr_o_16_, data_addr_o_15_, data_addr_o_14_, data_addr_o_13_, data_addr_o_12_, data_addr_o_11_, data_addr_o_10_, data_addr_o_9_, data_addr_o_8_, data_addr_o_7_, data_addr_o_6_, data_addr_o_5_, data_addr_o_4_, data_addr_o_3_, data_addr_o_2_, data_wdata_o_31_, data_wdata_o_30_, data_wdata_o_29_, data_wdata_o_28_, data_wdata_o_27_, data_wdata_o_26_, data_wdata_o_25_, data_wdata_o_24_, data_wdata_o_23_, data_wdata_o_22_, data_wdata_o_21_, data_wdata_o_20_, data_wdata_o_19_, data_wdata_o_18_, data_wdata_o_17_, data_wdata_o_16_, data_wdata_o_15_, data_wdata_o_14_, data_wdata_o_13_, data_wdata_o_12_, data_wdata_o_11_, data_wdata_o_10_, data_wdata_o_9_, data_wdata_o_8_, data_wdata_o_7_, data_wdata_o_6_, data_wdata_o_5_, data_wdata_o_4_, data_wdata_o_3_, data_wdata_o_2_, data_wdata_o_1_, data_wdata_o_0_, rf_we_wb_o, rf_wdata_wb_ecc_o_31_, rf_wdata_wb_ecc_o_30_, rf_wdata_wb_ecc_o_29_, rf_wdata_wb_ecc_o_28_, rf_wdata_wb_ecc_o_27_, rf_wdata_wb_ecc_o_26_, rf_wdata_wb_ecc_o_25_, rf_wdata_wb_ecc_o_24_, rf_wdata_wb_ecc_o_23_, rf_wdata_wb_ecc_o_22_, rf_wdata_wb_ecc_o_21_, rf_wdata_wb_ecc_o_20_, rf_wdata_wb_ecc_o_19_, rf_wdata_wb_ecc_o_18_, rf_wdata_wb_ecc_o_17_, rf_wdata_wb_ecc_o_16_, rf_wdata_wb_ecc_o_15_, rf_wdata_wb_ecc_o_14_, rf_wdata_wb_ecc_o_13_, rf_wdata_wb_ecc_o_12_, rf_wdata_wb_ecc_o_11_, rf_wdata_wb_ecc_o_10_, rf_wdata_wb_ecc_o_9_, rf_wdata_wb_ecc_o_8_, rf_wdata_wb_ecc_o_7_, rf_wdata_wb_ecc_o_6_, rf_wdata_wb_ecc_o_5_, rf_wdata_wb_ecc_o_4_, rf_wdata_wb_ecc_o_3_, rf_wdata_wb_ecc_o_2_, rf_wdata_wb_ecc_o_1_, rf_wdata_wb_ecc_o_0_, irq_pending_o, core_busy_o, n14858, n15022, n15310, n15145, n15259, n14806, n15044, n15194, n15165, n15578, n15102, n15419, n14828, n15752, n15049, n14962, n15305, n15553, n14984, n14994, n15075, n15337, n14889, n15120, n15333, n15656, n14981, n15146, n15642, n15085, n15089, n15162, n15300, n15711, n15453, n14867, n15359, n15696, n14955, n15101, n14844, n14997, n15313, n15495, n15598, n15076, n14813, n14894, n15509, n15096, n15543, n15549, n15732, n15399, n15540, n14810, n15209, n15647, n15702, n15555, n14931, n15295, n15195, n15319, n15452, n15173, n15779, n15363, n15500, n14795, n14912, n15180, n15528, n15311, n15216, n15439, n15464, n15105, n15427, n15738, n15035, n15286, n15742, n15253, n14939, n15348, n15535, n15449, n15245, n15671, n15255, n15139, n15274, n15579, n15434, n15352, n15334, n15007, n14978, n15715, n15230, n15457, n14857, n14871, n15095, n15005, n15367, n15382, n15210, n15402, n15629, n15126, n15001, n14824, n15289, n15624, n15615, n15755, n15753, n15197, n15583, n15408, n14869, n15386, n15155, n15531, n14950, n14959, n15090, n14907, n15061, n15567, n15584, n15680, n15377, n14974, n15364, n15397, n15657, n15706, n15610, n14905, n14996, n15028, n14930, n14964, n15018, n15002, n15666, n15699, n15083, n15281, n15082, n15136, n15390, n15396, n15668, n15144, n15569, n15237, n15485, n15737, n15762, n14802, n15107, n15674, n15203, n14926, n15700, n15128, n15763, n15443, n15631, n14929, n15678, n14899, n14911, n15006, n15284, n15297, n15694, n14918, n15264, n15244, n14897, n15034, n15338, n15053, n15117, n14881, n15213, n15123, n14944, n14975, n14801, n15461, n15356, n15030, n15058, n15436, n15703, n14972, n15276, n14812, n15529, n15676, n15254, n15488, n15565, n15079, n15772, n15635, n15458, n15133, n14993, n15198, n15234, n15783, n14831, n14854, n15070, n15186, n15669, n14841, n15655, n14816, n15721, n15777, n15008, n15009, n15039, n15534, n15438, n15557, n15329, n15292, n15603, n15758, n15645, n15560, n15100, n15731, n15767, n15004, n15068, n15059, n15243, n14951, n14830, n14794, n14901, n15369, n15116, n14970, n15413, n15526, n15476, n15091, n14792, n15312, n15403, n20894, n14935, n15564, n14922, n15723, n14908, n15539, n15612, n15520, n14868, n15507, n15024, n15094, n15646, n15071, n15472, n15287, n15012, n14875, n15092, n15221, n15261, n14878, n14843, n15063, n15505, n15527, n14840, n15684, n14838, n14865, n15681, n15558, n15391, n15351, n15563, n15045, n15097, n15229, n15317, n14800, n14803, n15484, n15219, n15185, n14882, n14827, n15335, n15459, n15513, n14913, n15157, n15478, n15545, n15099, n15160, n15395, n15316, n15379, n14851, n15775, n15542, n15613, n15191, n14872, n15582, n15764, n14988, n15704, n15770, n14823, n14814, n15471, n14817, n15376, n15258, n15052, n15639, n15765, n15291, n14876, n15188, n14917, n15381, n15416, n15087, n15371, n14808, n15062, n15538, n15698, n14958, n14826, n15228, n15760, n15013, n15246, n15130, n14973, n15385, n15410, n15027, n15415, n15514, n15278, n15033, n15400, n15423, n15517, n15345, n15301, n15781, n14825, n14921, n15113, n15304, n15622, n15620, n15486, n15498, n14938, n15588, n15277, n15242, n14864, n15283, n15321, n14859, n15177, n15554, n14885, n15435, n15648, n15153, n15709, n15282, n15437, n14999, n14799, n15467, n15548, n14804, n15241, n15720, n15134, n15406, n15456, n15586, n15651, n15688, n15362, n15743, n14797, n15215, n15633, n15510, n15019, n15572, n15341, n14880, n15773, n15469, n14989, n14998, n15183, n14941, n15078, n14822, n15148, n14942, n14990, n15468, n15129, n15235, n15477, n15734, n15231, n15710, n15636, n15201, n15626, n15315, n15728, n15644, n15273, n15205, n15239, n15298, n15294, n15414, n15649, n14874, n15643, n15675, n15025, n15733, n15374, n15713, n15494, n15223, n15663, n15550, n15530, n15673, n14916, n15288, n15296, n15330, n15121, n14957, n15141, n15306, n15614, n15693, n15716, n15761, n14956, n15735, n15232, n15200, n15060, n15571, n14960, n15621, n15072, n15174, n15451, n15159, n14818, n15618, n14948, n14850, n15346, n14952, n15503, n15279, n15178, n14967, n15522, n15263, n15533, n14963, n14842, n15041, n15577, n14992, n15506, n14853, n15780, n14852, n15236, n15532, n15428, n15179, n15418, n15450, n15115, n14979, n15591, n15354, n14886, n14892, n15623, n15559, n14968, n15320, n15175, n15525, n15653, n15110, n15192, n14919, n14821, n15574, n14947, n15048, n15014, n15168, n15344, n14811, n15054, n15166, n15260, n15608, n15508, n15405, n14820, n14928, n15566, n14903, n14891, n15616, n15147, n15524, n14927, n15073, n14923, n15328, n15609, n15705, n15782, n14914, n15055, n15754, n14896, n15679, n15164, n15086, n15501, n14848, n15124, n15685, n15491, n15015, n15140, n15360, n15474, n15740, n14796, n15190, n15447, n15098, n14870, n14977, n15302, n15023, n14982, n15046, n15339, n15718, n15430, n14835, n15189, n15251, n15778, n15383, n15003, n15431, n15512, n15275, n15463, n15421, n15519, n15161, n15355, n15561, n15208, n14863, n15714, n15749, n15759, n15632, n15365, n15747, n14860, n15156, n15187, n15604, n15336, n15375, n15342, n15404, n15257, n15118, n15499, n15585, n15575, n15619, n15163, n15701, n15465, n15167, n15268, n15370, n15487, n15220, n15088, n15309, n15521, n15625, n14845, n14856, n14887, n15067, n15470, n15768, n15171, n15446, n15248, n15687, n15412, n15043, n15104, n14890, n14936, n15247, n14991, n15384, n15690, n14834, n15717, n14966, n15448, n15432, n15659, n15686, n15212, n15020, n15303, n15214, n15314, n15181, n15047, n15154, n15401, n14862, n14980, n15318, n15589, n14924, n15462, n15016, n14940, n15358, n15409, n14829, n14920, n15712, n15460, n14866, n15143, n14832, n14855, n15466, n14847, n15056, n15637, n15660, n15597, n15125, n14805, n15069, n15581, n15724, n15211, n15222, n15066, n15176, n15592, n15158, n15373, n15601, n15748, n14888, n15587, n15349, n15350, n14949, n14971, n15372, n15599, n14983, n15347, n15380, n15650, n15727, n14877, n15325, n15324, n15119, n15106, n15407, n15233, n15691, n14833, n15745, n15327, n14986, n15425, n15149, n15602, n15692, n15658, n15207, n14807, n15594, n15766, n14879, n15111, n15475, n15152, n15299, n14965, n15455, n15667, n15093, n15326, n15249, n15074, n15661, n15473, n15172, n15388, n15000, n15227, n15114, n15366, n15307, n15689, n14861, n15638, n15184, n15593, n14809, n15280, n15017, n14849, n15193, n14987, n15265, n14898, n14925, n15109, n15011, n15270, n15562, n15739, n15196, n15708, n14895, n15741, n15677, n15670, n15672, n15323, n15511, n15695, n15361, n15537, n15634, n15081, n15202, n15256, n15750, n15084, n15343, n15262, n15454, n15568, n14904, n15142, n14946, n15627, n15040, n15744, n15445, n14793, n15151, n15077, n15132, n15544, n15665, n14883, n15080, n15226, n15492, n14839, n15523, n15417, n15387, n15206, n15641, n14976, n15150, n15607, n15751, n15340, n14954, n15444, n15021, n15285, n15757, n15774, n15331, n15037, n15240, n15730, n15489, n15722, n15606, n15010, n15424, n15547, n15392, n15064, n15138, n14884, n15199, n15411, n15652, n15576, n15429, n14943, n15029, n14934, n15269, n15422, n14969, n14900, n15218, n15332, n14798, n15137, n15042, n14995, n15420, n15122, n15182, n15490, n14873, n15169, n14915, n15515, n15611, n15725, n14910, n15031, n15026, n15573, n15493, n15496, n15719, n14893, n15112, n15252, n15426, n15127, n15536, n15441, n15541, n15204, n15442, n15271, n14906, n15483, n15580, n14937, n15596, n15225, n15726, n15038, n15065, n15697, n15481, n15497, n15518, n15736, n15272, n14815, n14902, n15398, n15322, n15353, n15546, n15502, n14945, n15504, n15050, n15654, n15769, n15357, n15482, n15368, n14846, n15433, n15378, n14836, n15057, n15682, n14909, n15516, n15266, n15628, n15393, n15308, n15590, n15103, n14933, n15394, n20877, n15479, n15480, n15108, n15217, n15776, n15707, n15662, n15051, n15224, n15756, n14932, n14985, n15600, n15595, n15250, n15389, n15640, n14953, n15729, n15551, n15440, n15552, n14961, n15238, n15605, n15135, n15630, n15664, n15570, n15746, n14819, n15267, n15290, n15683, n14837, n15032, n15170, n15771, n15036, n15131, n15293, n15617;
wire if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N38, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N37, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N36, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N35, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N34, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N33, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N32, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N31, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N30, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N29, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N28, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N27, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N26, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N25, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N24, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N23, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N22, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N21, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N20, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N19, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N18, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N17, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N16, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N15, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N14, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N13, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N12, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N11, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N9, id_stage_i_controller_i_N288, id_stage_i_controller_i_N287, id_stage_i_controller_i_N286, id_stage_i_controller_i_N285, id_stage_i_controller_i_N284, id_stage_i_controller_i_N283, id_stage_i_controller_i_N282, id_stage_i_controller_i_N281, id_stage_i_controller_i_N280, id_stage_i_controller_i_N279, id_stage_i_controller_i_N278, id_stage_i_controller_i_N277, id_stage_i_controller_i_N276, id_stage_i_controller_i_N275, id_stage_i_controller_i_N274, id_stage_i_controller_i_N273, id_stage_i_controller_i_N272, id_stage_i_controller_i_N271, id_stage_i_controller_i_N270, id_stage_i_controller_i_N269, id_stage_i_controller_i_N268, id_stage_i_controller_i_N267, id_stage_i_controller_i_N266, id_stage_i_controller_i_N265, id_stage_i_controller_i_N264, id_stage_i_controller_i_N263, id_stage_i_controller_i_N262, id_stage_i_controller_i_N261, id_stage_i_controller_i_N260, id_stage_i_controller_i_N259, id_stage_i_controller_i_N258, ex_block_i_alu_is_equal_result, ex_block_i_alu_i_N294, ex_block_i_gen_multdiv_fast_multdiv_i_N221, ex_block_i_gen_multdiv_fast_multdiv_i_N220, ex_block_i_gen_multdiv_fast_multdiv_i_N219, ex_block_i_gen_multdiv_fast_multdiv_i_N218, ex_block_i_gen_multdiv_fast_multdiv_i_sign_b, ex_block_i_gen_multdiv_fast_multdiv_i_sign_a, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N68, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N67, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N66, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N65, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N64, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N63, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N62, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N61, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N60, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N59, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N58, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N57, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N56, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N55, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N54, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N53, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N52, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N51, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N50, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N49, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N48, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N47, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N46, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N45, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N44, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N43, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N42, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N41, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N40, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N39, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N38, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N37, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N36, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N35, n32, n33, n34, n35, n36, n37, n38, n39, n42, n43, n44, n45, n47, n48, n49, n50, n51, n52, n54, n55, n56, n58, n59, n60, n61, n65, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81, n83, n85, n86, n87, n88, n89, n90, n92, n94, n95, n96, n97, n98, n99, n101, n102, n104, n105, n106, n107, n108, n109, n110, n111, n113, n114, n115, n116, n117, n118, n119, n120, n121, n123, n124, n125, n126, n127, n128, n129, n131, n132, n133, n134, n137, n138, n139, n140, n141, n142, n144, n145, n146, n147, n148, n149, n150, n151, n154, n156, n157, n158, n159, n160, n161, n162, n163, n165, n166, n169, n170, n171, n172, n173, n174, n175, n176, n177, n179, n180, n181, n182, n185, n186, n187, n188, n189, n190, n192, n193, n194, n195, n196, n197, n198, n199, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n213, n214, n215, n216, n217, n218, n219, n220, n222, n223, n224, n225, n228, n229, n230, n231, n232, n233, n235, n236, n237, n238, n239, n240, n241, n242, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n264, n265, n266, n267, n270, n271, n272, n273, n274, n275, n277, n278, n279, n280, n281, n282, n283, n284, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n305, n306, n307, n308, n311, n312, n313, n314, n315, n316, n318, n319, n320, n321, n322, n323, n324, n325, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n346, n347, n348, n349, n352, n353, n354, n355, n356, n357, n359, n360, n361, n363, n365, n366, n367, n368, n370, n371, n373, n374, n376, n378, n379, n380, n381, n382, n383, n384, n385, n386, n388, n389, n390, n391, n394, n395, n399, n400, n401, n402, n403, n404, n405, n406, n409, n410, n411, n412, n413, n414, n415, n416, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n431, n432, n433, n434, n436, n437, n440, n441, n442, n443, n444, n445, n447, n448, n449, n450, n451, n452, n453, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n468, n469, n470, n471, n472, n473, n474, n476, n477, n478, n479, n482, n483, n484, n485, n486, n487, n488, n489, n492, n493, n494, n495, n496, n497, n498, n499, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n514, n515, n516, n517, n519, n520, n522, n523, n524, n525, n526, n527, n528, n529, n532, n533, n534, n535, n536, n537, n538, n539, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n554, n555, n556, n557, n559, n560, n562, n563, n564, n565, n566, n567, n568, n569, n572, n573, n574, n575, n576, n577, n578, n579, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n594, n595, n596, n597, n599, n600, n602, n603, n604, n605, n606, n607, n608, n609, n612, n613, n614, n615, n616, n617, n618, n619, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n634, n635, n636, n637, n639, n640, n642, n643, n644, n645, n646, n647, n648, n649, n652, n653, n654, n655, n656, n657, n658, n659, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n673, n674, n675, n676, n677, n678, n680, n681, n682, n683, n684, n685, n686, n687, n690, n691, n692, n693, n694, n695, n696, n697, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n711, n712, n713, n714, n715, n716, n718, n719, n720, n721, n722, n723, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n748, n749, n750, n751, n752, n753, n755, n756, n757, n758, n759, n760, n762, n763, n765, n766, n767, n768, n769, n770, n771, n772, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n786, n787, n788, n789, n790, n791, n793, n794, n795, n796, n797, n798, n800, n801, n803, n804, n805, n806, n807, n808, n809, n810, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n824, n825, n826, n827, n828, n829, n832, n833, n834, n835, n836, n837, n839, n840, n842, n843, n844, n845, n846, n847, n848, n849, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n863, n864, n865, n866, n867, n868, n871, n872, n873, n874, n875, n876, n878, n879, n880, n881, n882, n883, n884, n885, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n913, n914, n915, n916, n917, n918, n920, n921, n923, n924, n925, n926, n927, n928, n929, n930, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n944, n945, n946, n947, n948, n949, n952, n953, n954, n955, n956, n957, n959, n960, n962, n963, n964, n965, n966, n967, n968, n969, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n983, n984, n985, n986, n987, n988, n991, n992, n993, n994, n995, n996, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1021, n1022, n1023, n1024, n1025, n1026, n1029, n1030, n1031, n1032, n1033, n1034, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1048, n1049, n1050, n1051, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1063, n1064, n1065, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1079, n1080, n1081, n1082, n1084, n1085, n1088, n1089, n1090, n1091, n1092, n1093, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1127, n1128, n1129, n1130, n1131, n1132, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1166, n1167, n1168, n1169, n1170, n1171, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1205, n1206, n1207, n1208, n1209, n1210, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1244, n1245, n1246, n1247, n1248, n1249, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1283, n1284, n1285, n1286, n1287, n1288, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1311, n1312, n1313, n1314, n1315, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1362, n1363, n1364, n1365, n1366, n1368, n1372, n1373, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1401, n1404, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1415, n1416, n1417, n1418, n1419, n1420, n1422, n1423, n1426, n1427, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1442, n1443, n1444, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1504, n1505, n1507, n1508, n1509, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1520, n1521, n1522, n1524, n1525, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1536, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1558, n1559, n1560, n1561, n1562, n1564, n1565, n1566, n1567, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1606, n1607, n1608, n1610, n1611, n1613, n1614, n1616, n1617, n1619, n1620, n1622, n1623, n1625, n1626, n1628, n1629, n1631, n1632, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1653, n1654, n1655, n1656, n1657, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1670, n1671, n1673, n1674, n1676, n1677, n1679, n1680, n1682, n1683, n1685, n1686, n1687, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1698, n1699, n1700, n1701, n1704, n1705, n1706, n1708, n1709, n1710, n1712, n1713, n1715, n1716, n1718, n1719, n1721, n1722, n1724, n1725, n1727, n1728, n1730, n1731, n1733, n1734, n1736, n1737, n1739, n1740, n1742, n1743, n1745, n1746, n1748, n1749, n1751, n1752, n1754, n1755, n1757, n1758, n1760, n1761, n1763, n1764, n1766, n1767, n1769, n1770, n1772, n1773, n1775, n1776, n1778, n1779, n1781, n1782, n1784, n1785, n1787, n1788, n1790, n1791, n1793, n1794, n1796, n1797, n1799, n1800, n1802, n1803, n1805, n1806, n1808, n1809, n1811, n1812, n1814, n1815, n1817, n1818, n1820, n1821, n1823, n1824, n1826, n1827, n1829, n1830, n1832, n1833, n1835, n1836, n1838, n1839, n1841, n1842, n1844, n1845, n1847, n1848, n1850, n1851, n1853, n1854, n1856, n1857, n1859, n1860, n1862, n1863, n1865, n1866, n1868, n1869, n1871, n1872, n1874, n1875, n1877, n1878, n1880, n1881, n1883, n1884, n1885, n1889, n1890, n1893, n1894, n1897, n1898, n1901, n1902, n1904, n1905, n1907, n1908, n1910, n1911, n1913, n1914, n1916, n1917, n1919, n1920, n1923, n1924, n1927, n1928, n1931, n1932, n1935, n1936, n1939, n1940, n1943, n1944, n1947, n1948, n1951, n1952, n1954, n1955, n1958, n1959, n1961, n1962, n1965, n1966, n1969, n1970, n1973, n1974, n1977, n1978, n1981, n1982, n1985, n1986, n1989, n1990, n1993, n1994, n1996, n1997, n2000, n2001, n2003, n2004, n2005, n2006, n2007, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2018, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2053, n2054, n2055, n2056, n2058, n2059, n2060, n2061, n2062, n2064, n2065, n2066, n2067, n2068, n2069, n2071, n2072, n2074, n2075, n2077, n2078, n2080, n2081, n2082, n2084, n2085, n2087, n2088, n2090, n2091, n2093, n2094, n2096, n2097, n2098, n2099, n2100, n2102, n2103, n2104, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2125, n2126, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2152, n2154, n2155, n2156, n2157, n2159, n2160, n2161, n2162, n2163, n2164, n2166, n2167, n2168, n2169, n2170, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2197, n2198, n2199, n2202, n2203, n2204, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2214, n2215, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2229, n2230, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2245, n2246, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2258, n2259, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2279, n2280, n2281, n2282, n2283, n2284, n2286, n2287, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2302, n2303, n2304, n2305, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2315, n2316, n2318, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2329, n2330, n2332, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2351, n2352, n2354, n2355, n2356, n2358, n2359, n2360, n2361, n2363, n2365, n2366, n2367, n2368, n2370, n2371, n2373, n2374, n2375, n2376, n2377, n2378, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2412, n2413, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2468, n2470, n2471, n2472, n2474, n2475, n2476, n2477, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2489, n2491, n2492, n2494, n2495, n2496, n2497, n2498, n2500, n2501, n2503, n2504, n2505, n2508, n2509, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2560, n2561, n2562, n2563, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2578, n2579, n2581, n2582, n2584, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2607, n2608, n2610, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2635, n2636, n2638, n2639, n2640, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2673, n2674, n2675, n2676, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2689, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2704, n2705, n2707, n2708, n2709, n2710, n2711, n2712, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2794, n2795, n2797, n2798, n2799, n2800, n2801, n2803, n2804, n2806, n2807, n2808, n2809, n2811, n2812, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2830, n2831, n2832, n2833, n2835, n2836, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2876, n2877, n2879, n2880, n2881, n2882, n2884, n2885, n2887, n2888, n2889, n2890, n2892, n2893, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3024, n3025, n3027, n3028, n3029, n3030, n3032, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3045, n3047, n3048, n3049, n3050, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3356, n3357, n3358, n3359, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3500, n3501, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3611, n3612, n3613, n3615, n3616, n3618, n3619, n3621, n3622, n3624, n3625, n3627, n3628, n3630, n3631, n3633, n3634, n3636, n3637, n3639, n3640, n3642, n3643, n3645, n3646, n3648, n3649, n3651, n3652, n3654, n3655, n3657, n3658, n3660, n3661, n3663, n3664, n3666, n3667, n3669, n3670, n3672, n3673, n3675, n3676, n3678, n3679, n3681, n3682, n3684, n3685, n3687, n3688, n3690, n3691, n3693, n3694, n3696, n3697, n3699, n3700, n3702, n3703, n3704, n3705, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4004, n4005, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4054, n4056, n4057, n4058, n4059, n4060, n4061, n4063, n4064, n4066, n4067, n4068, n4069, n4071, n4072, n4074, n4075, n4077, n4078, n4080, n4081, n4083, n4084, n4086, n4087, n4089, n4090, n4092, n4093, n4095, n4096, n4098, n4099, n4101, n4102, n4104, n4105, n4107, n4108, n4110, n4111, n4113, n4114, n4116, n4117, n4119, n4120, n4122, n4123, n4125, n4126, n4128, n4129, n4131, n4132, n4134, n4135, n4137, n4138, n4140, n4141, n4143, n4144, n4146, n4147, n4149, n4150, n4152, n4153, n4155, n4156, n4158, n4159, n4161, n4162, n4164, n4165, n4167, n4168, n4170, n4171, n4173, n4174, n4176, n4177, n4179, n4180, n4182, n4183, n4185, n4186, n4188, n4189, n4191, n4192, n4194, n4195, n4197, n4198, n4200, n4201, n4203, n4204, n4206, n4207, n4209, n4210, n4212, n4213, n4215, n4216, n4218, n4219, n4221, n4222, n4224, n4225, n4227, n4228, n4230, n4231, n4233, n4234, n4236, n4237, n4239, n4240, n4242, n4243, n4245, n4246, n4248, n4249, n4253, n4254, n4256, n4257, n4258, n4260, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4270, n4271, n4272, n4273, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4285, n4286, n4287, n4288, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4308, n4309, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4327, n4328, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4346, n4347, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4365, n4366, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4384, n4385, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4403, n4404, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4420, n4421, n4422, n4423, n4425, n4426, n4427, n4428, n4430, n4431, n4432, n4433, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4443, n4444, n4445, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4457, n4458, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4478, n4479, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4497, n4498, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4518, n4519, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4539, n4540, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4560, n4561, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4581, n4582, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4602, n4603, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4623, n4624, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4644, n4645, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4665, n4666, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4686, n4687, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4707, n4708, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4746, n4747, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4767, n4768, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4788, n4789, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4810, n4811, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4829, n4830, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4848, n4849, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4867, n4868, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4886, n4887, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4905, n4906, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4929, n4930, n4932, n4933, n4934, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4952, n4953, n4955, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4970, n4972, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4994, n4995, n4996, n4998, n5000, n5001, n5002, n5003, n5004, n5005, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5022, n5023, n5026, n5027, n5028, n5029, n5030, n5031, n5033, n5035, n5036, n5037, n5038, n5039, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5072, n5073, n5074, n5075, n5077, n5078, n5079, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5112, n5113, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5159, n5160, n5161, n5162, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5180, n5182, n5183, n5184, n5185, n5186, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5196, n5197, n5198, n5200, n5201, n5202, n5204, n5205, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5232, n5233, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5253, n5254, n5255, n5256, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5266, n5267, n5268, n5269, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5280, n5281, n5283, n5284, n5286, n5287, n5289, n5290, n5292, n5293, n5295, n5296, n5298, n5299, n5301, n5302, n5304, n5305, n5307, n5308, n5310, n5311, n5313, n5314, n5316, n5317, n5319, n5320, n5322, n5323, n5325, n5326, n5328, n5329, n5331, n5332, n5334, n5335, n5337, n5338, n5340, n5341, n5343, n5344, n5346, n5347, n5349, n5350, n5352, n5353, n5355, n5356, n5358, n5359, n5361, n5362, n5364, n5365, n5367, n5368, n5370, n5371, n5372, n5374, n5375, n5376, n5377, n5378, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5390, n5391, n5392, n5393, n5395, n5396, n5397, n5398, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5426, n5427, n5428, n5429, n5431, n5432, n5433, n5434, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5478, n5479, n5480, n5481, n5483, n5484, n5485, n5486, n5488, n5489, n5490, n5491, n5493, n5494, n5495, n5496, n5498, n5499, n5500, n5501, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5516, n5517, n5518, n5519, n5521, n5522, n5523, n5524, n5526, n5527, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5559, n5560, n5562, n5566, n5567, n5569, n5571, n5573, n5574, n5575, n5578, n5579, n5580, n5581, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5690, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5818, n5820, n5821, n5822, n5823, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6183, n6184, n6185, n6186, n6187, n6188, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6517, n6518, n6519, n6520, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6545, n6546, n6547, n6549, n6550, n6552, n6554, n6555, n6556, n6557, n6558, n6561, n6562, n6563, n6564, n6565, n6568, n6569, n6570, n6571, n6574, n6575, n6576, n6577, n6580, n6581, n6582, n6583, n6586, n6587, n6588, n6589, n6592, n6593, n6594, n6595, n6598, n6599, n6600, n6601, n6604, n6605, n6606, n6607, n6610, n6611, n6612, n6613, n6616, n6617, n6618, n6619, n6622, n6623, n6624, n6625, n6628, n6629, n6630, n6631, n6634, n6635, n6636, n6637, n6640, n6641, n6642, n6643, n6646, n6647, n6648, n6649, n6652, n6653, n6654, n6655, n6658, n6659, n6660, n6661, n6664, n6665, n6666, n6667, n6670, n6671, n6672, n6673, n6676, n6677, n6678, n6679, n6682, n6683, n6684, n6685, n6688, n6689, n6690, n6691, n6694, n6695, n6697, n6698, n6699, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6813, n6814, n6815, n6816, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7059, n7060, n7061, n7062, n7063, n7064, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7074, n7075, n7076, n7077, n7078, n7081, n7082, n7084, n7107, n7108, n7109, n7110, n7113, n7114, n7123, n7124, n7133, n7134, n7143, n7144, n7147, n7148, n7150, n7151, n7156, n7157, n7160, n7161, n7164, n7165, n7167, n7168, n7170, n7171, n7173, n7174, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7255, n7256, n7257, n7260, n7261, n7263, n7264, n7266, n7267, n7269, n7270, n7272, n7273, n7275, n7276, n7278, n7279, n7281, n7282, n7284, n7285, n7287, n7288, n7289, n7290, n7292, n7293, n7295, n7296, n7298, n7299, n7301, n7302, n7304, n7305, n7307, n7308, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7601, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7649, n7650, n7651, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7683, n7684, n7685, n7686, n7687, n7688, n7690, n7691, n7692, n7693, n7694, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7704, n7705, n7707, n7708, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7728, n7729, n7730, n7731, n7732, n7733, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7780, n7781, n7783, n7784, n7786, n7787, n7788, n7789, n7790, n7791, n7793, n7794, n7795, n7796, n7797, n7799, n7800, n7801, n7802, n7803, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7862, n7863, n7864, n7865, n7867, n7868, n7869, n7870, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8056, n8057, n8058, n8060, n8061, n8062, n8063, n8065, n8068, n8069, n8070, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8091, n8092, n8093, n8094, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8106, n8107, n8108, n8111, n8112, n8113, n8115, n8116, n8117, n8118, n8119, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8308, n8309, n8310, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8424, n8426, n8429, n8430, n8431, n8432, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8565, n8566, n8567, n8568, n8569, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8595, n8596, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8885, n8886, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9843, n9844, n9845, n9846, n9848, n9849, n9850, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9911, n9912, n9913, n9914, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9944, n9945, n9947, n9948, n9949, n9950, n9952, n9953, n9954, n9955, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10156, n10157, n10158, n10159, n10160, n10161, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10182, n10183, n10184, n10185, n10187, n10188, n10189, n10191, n10192, n10193, n10196, n10197, n10198, n10199, n10201, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10295, n10296, n10297, n10298, n10300, n10301, n10302, n10303, n10304, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10403, n10404, n10405, n10406, n10407, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10431, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10444, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_15_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_16_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_17_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_18_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_19_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_20_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_21_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_22_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_23_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_24_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_25_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_26_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_27_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_28_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_29_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_30_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_31_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_15_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_16_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_17_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_18_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_19_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_20_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_21_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_22_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_23_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_24_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_25_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_26_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_27_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_28_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_29_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_30_, dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_31_, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fifo_i_add_146_B_1_, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_add_243_A_1_, n15794, n15795, n15796, n15797, n15801, n15802, n15808, n15811, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668, alu_operand_b_ex_4, alu_operand_b_ex_3, alu_operand_b_ex_2, alu_operand_b_ex_1, alu_adder_result_ex_1, alu_adder_result_ex_0, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_31, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_30, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_29, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_28, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_27, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_26, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_25, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_24, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_23, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_22, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_21, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_20, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_19, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_18, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_17, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_16, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_15, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_14, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_13, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_12, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_11, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_10, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_9, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_8, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_7, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_6, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_5, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_4, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_3, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_2, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_31, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_30, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_29, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_28, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_27, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_26, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_25, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_24, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_23, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_22, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_21, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_20, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_19, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_18, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_17, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_16, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_15, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_14, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_13, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_12, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_11, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_10, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_9, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_8, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_7, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_6, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_5, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_4, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_3, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_2, if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_1, ex_block_i_alu_i_shift_result_ext_signed_30, ex_block_i_alu_i_shift_result_ext_signed_29, ex_block_i_alu_i_shift_result_ext_signed_28, ex_block_i_alu_i_shift_result_ext_signed_27, ex_block_i_alu_i_shift_result_ext_signed_26, ex_block_i_alu_i_shift_result_ext_signed_25, ex_block_i_alu_i_shift_result_ext_signed_24, ex_block_i_alu_i_shift_result_ext_signed_23, ex_block_i_alu_i_shift_result_ext_signed_22, ex_block_i_alu_i_shift_result_ext_signed_21, ex_block_i_alu_i_shift_result_ext_signed_20, ex_block_i_alu_i_shift_result_ext_signed_19, ex_block_i_alu_i_shift_result_ext_signed_18, ex_block_i_alu_i_shift_result_ext_signed_17, ex_block_i_alu_i_shift_result_ext_signed_16, ex_block_i_alu_i_shift_operand_31, ex_block_i_alu_i_shift_operand_0, ex_block_i_alu_i_shift_amt_compl_4, ex_block_i_alu_i_shift_amt_compl_3, ex_block_i_alu_i_shift_amt_compl_2, ex_block_i_alu_i_shift_amt_compl_1, ex_block_i_alu_i_shift_amt_compl_0, ex_block_i_alu_i_shift_amt_4, ex_block_i_alu_i_shift_amt_3, ex_block_i_alu_i_shift_amt_2, ex_block_i_alu_i_shift_amt_1, ex_block_i_alu_i_shift_amt_0, ex_block_i_alu_i_adder_in_b_32, ex_block_i_alu_i_adder_in_b_31, ex_block_i_alu_i_adder_in_b_30, ex_block_i_alu_i_adder_in_b_29, ex_block_i_alu_i_adder_in_b_28, ex_block_i_alu_i_adder_in_b_27, ex_block_i_alu_i_adder_in_b_26, ex_block_i_alu_i_adder_in_b_25, ex_block_i_alu_i_adder_in_b_24, ex_block_i_alu_i_adder_in_b_23, ex_block_i_alu_i_adder_in_b_22, ex_block_i_alu_i_adder_in_b_21, ex_block_i_alu_i_adder_in_b_20, ex_block_i_alu_i_adder_in_b_19, ex_block_i_alu_i_adder_in_b_18, ex_block_i_alu_i_adder_in_b_17, ex_block_i_alu_i_adder_in_b_16, ex_block_i_alu_i_adder_in_b_15, ex_block_i_alu_i_adder_in_b_14, ex_block_i_alu_i_adder_in_b_13, ex_block_i_alu_i_adder_in_b_12, ex_block_i_alu_i_adder_in_b_11, ex_block_i_alu_i_adder_in_b_10, ex_block_i_alu_i_adder_in_b_9, ex_block_i_alu_i_adder_in_b_8, ex_block_i_alu_i_adder_in_b_7, ex_block_i_alu_i_adder_in_b_6, ex_block_i_alu_i_adder_in_b_5, ex_block_i_alu_i_adder_in_b_4, ex_block_i_alu_i_adder_in_b_3, ex_block_i_alu_i_adder_in_b_2, ex_block_i_alu_i_adder_in_b_1, ex_block_i_alu_i_adder_in_a_31, ex_block_i_alu_i_adder_in_a_30, ex_block_i_alu_i_adder_in_a_29, ex_block_i_alu_i_adder_in_a_28, ex_block_i_alu_i_adder_in_a_27, ex_block_i_alu_i_adder_in_a_26, ex_block_i_alu_i_adder_in_a_25, ex_block_i_alu_i_adder_in_a_24, ex_block_i_alu_i_adder_in_a_23, ex_block_i_alu_i_adder_in_a_22, ex_block_i_alu_i_adder_in_a_21, ex_block_i_alu_i_adder_in_a_20, ex_block_i_alu_i_adder_in_a_19, ex_block_i_alu_i_adder_in_a_18, ex_block_i_alu_i_adder_in_a_17, ex_block_i_alu_i_adder_in_a_16, ex_block_i_alu_i_adder_in_a_15, ex_block_i_alu_i_adder_in_a_14, ex_block_i_alu_i_adder_in_a_13, ex_block_i_alu_i_adder_in_a_12, ex_block_i_alu_i_adder_in_a_11, ex_block_i_alu_i_adder_in_a_10, ex_block_i_alu_i_adder_in_a_9, ex_block_i_alu_i_adder_in_a_8, ex_block_i_alu_i_adder_in_a_7, ex_block_i_alu_i_adder_in_a_6, ex_block_i_alu_i_adder_in_a_5, ex_block_i_alu_i_adder_in_a_4, ex_block_i_alu_i_adder_in_a_3, ex_block_i_alu_i_adder_in_a_2, ex_block_i_alu_i_adder_in_a_1, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_31, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_30, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_29, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_28, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_27, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_26, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_25, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_24, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_23, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_22, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_21, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_20, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_19, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_18, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_17, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_16, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_15, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_14, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_13, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_12, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_11, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_10, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_9, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_8, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_7, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_6, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_5, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_4, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_3, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_2, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_1, ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_0, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_33, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_32, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_31, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_30, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_29, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_28, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_27, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_26, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_25, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_24, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_23, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_22, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_21, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_20, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_19, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_18, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_17, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_16, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_15, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_14, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_13, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_12, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_11, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_10, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_9, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_8, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_7, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_6, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_5, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_4, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_3, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_2, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_1, ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_0, ex_block_i_gen_multdiv_fast_multdiv_i_accum_33, ex_block_i_gen_multdiv_fast_multdiv_i_accum_32, ex_block_i_gen_multdiv_fast_multdiv_i_accum_31, ex_block_i_gen_multdiv_fast_multdiv_i_accum_30, ex_block_i_gen_multdiv_fast_multdiv_i_accum_29, ex_block_i_gen_multdiv_fast_multdiv_i_accum_28, ex_block_i_gen_multdiv_fast_multdiv_i_accum_27, ex_block_i_gen_multdiv_fast_multdiv_i_accum_26, ex_block_i_gen_multdiv_fast_multdiv_i_accum_25, ex_block_i_gen_multdiv_fast_multdiv_i_accum_24, ex_block_i_gen_multdiv_fast_multdiv_i_accum_23, ex_block_i_gen_multdiv_fast_multdiv_i_accum_22, ex_block_i_gen_multdiv_fast_multdiv_i_accum_21, ex_block_i_gen_multdiv_fast_multdiv_i_accum_20, ex_block_i_gen_multdiv_fast_multdiv_i_accum_19, ex_block_i_gen_multdiv_fast_multdiv_i_accum_18, ex_block_i_gen_multdiv_fast_multdiv_i_accum_17, ex_block_i_gen_multdiv_fast_multdiv_i_accum_16, ex_block_i_gen_multdiv_fast_multdiv_i_accum_15, ex_block_i_gen_multdiv_fast_multdiv_i_accum_14, ex_block_i_gen_multdiv_fast_multdiv_i_accum_13, ex_block_i_gen_multdiv_fast_multdiv_i_accum_12, ex_block_i_gen_multdiv_fast_multdiv_i_accum_11, ex_block_i_gen_multdiv_fast_multdiv_i_accum_10, ex_block_i_gen_multdiv_fast_multdiv_i_accum_9, ex_block_i_gen_multdiv_fast_multdiv_i_accum_8, ex_block_i_gen_multdiv_fast_multdiv_i_accum_7, ex_block_i_gen_multdiv_fast_multdiv_i_accum_6, ex_block_i_gen_multdiv_fast_multdiv_i_accum_5, ex_block_i_gen_multdiv_fast_multdiv_i_accum_4, ex_block_i_gen_multdiv_fast_multdiv_i_accum_3, ex_block_i_gen_multdiv_fast_multdiv_i_accum_2, ex_block_i_gen_multdiv_fast_multdiv_i_accum_1, ex_block_i_gen_multdiv_fast_multdiv_i_accum_0, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_1, ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0, cs_registers_i_mcycle_counter_i_counter_upd_63, cs_registers_i_mcycle_counter_i_counter_upd_62, cs_registers_i_mcycle_counter_i_counter_upd_61, cs_registers_i_mcycle_counter_i_counter_upd_60, cs_registers_i_mcycle_counter_i_counter_upd_59, cs_registers_i_mcycle_counter_i_counter_upd_58, cs_registers_i_mcycle_counter_i_counter_upd_57, cs_registers_i_mcycle_counter_i_counter_upd_56, cs_registers_i_mcycle_counter_i_counter_upd_55, cs_registers_i_mcycle_counter_i_counter_upd_54, cs_registers_i_mcycle_counter_i_counter_upd_53, cs_registers_i_mcycle_counter_i_counter_upd_52, cs_registers_i_mcycle_counter_i_counter_upd_51, cs_registers_i_mcycle_counter_i_counter_upd_50, cs_registers_i_mcycle_counter_i_counter_upd_49, cs_registers_i_mcycle_counter_i_counter_upd_48, cs_registers_i_mcycle_counter_i_counter_upd_47, cs_registers_i_mcycle_counter_i_counter_upd_46, cs_registers_i_mcycle_counter_i_counter_upd_45, cs_registers_i_mcycle_counter_i_counter_upd_44, cs_registers_i_mcycle_counter_i_counter_upd_43, cs_registers_i_mcycle_counter_i_counter_upd_42, cs_registers_i_mcycle_counter_i_counter_upd_41, cs_registers_i_mcycle_counter_i_counter_upd_40, cs_registers_i_mcycle_counter_i_counter_upd_39, cs_registers_i_mcycle_counter_i_counter_upd_38, cs_registers_i_mcycle_counter_i_counter_upd_37, cs_registers_i_mcycle_counter_i_counter_upd_36, cs_registers_i_mcycle_counter_i_counter_upd_35, cs_registers_i_mcycle_counter_i_counter_upd_34, cs_registers_i_mcycle_counter_i_counter_upd_33, cs_registers_i_mcycle_counter_i_counter_upd_32, cs_registers_i_mcycle_counter_i_counter_upd_31, cs_registers_i_mcycle_counter_i_counter_upd_30, cs_registers_i_mcycle_counter_i_counter_upd_29, cs_registers_i_mcycle_counter_i_counter_upd_28, cs_registers_i_mcycle_counter_i_counter_upd_27, cs_registers_i_mcycle_counter_i_counter_upd_26, cs_registers_i_mcycle_counter_i_counter_upd_25, cs_registers_i_mcycle_counter_i_counter_upd_24, cs_registers_i_mcycle_counter_i_counter_upd_23, cs_registers_i_mcycle_counter_i_counter_upd_22, cs_registers_i_mcycle_counter_i_counter_upd_21, cs_registers_i_mcycle_counter_i_counter_upd_20, cs_registers_i_mcycle_counter_i_counter_upd_19, cs_registers_i_mcycle_counter_i_counter_upd_18, cs_registers_i_mcycle_counter_i_counter_upd_17, cs_registers_i_mcycle_counter_i_counter_upd_16, cs_registers_i_mcycle_counter_i_counter_upd_15, cs_registers_i_mcycle_counter_i_counter_upd_14, cs_registers_i_mcycle_counter_i_counter_upd_13, cs_registers_i_mcycle_counter_i_counter_upd_12, cs_registers_i_mcycle_counter_i_counter_upd_11, cs_registers_i_mcycle_counter_i_counter_upd_10, cs_registers_i_mcycle_counter_i_counter_upd_9, cs_registers_i_mcycle_counter_i_counter_upd_8, cs_registers_i_mcycle_counter_i_counter_upd_7, cs_registers_i_mcycle_counter_i_counter_upd_6, cs_registers_i_mcycle_counter_i_counter_upd_5, cs_registers_i_mcycle_counter_i_counter_upd_4, cs_registers_i_mcycle_counter_i_counter_upd_3, cs_registers_i_mcycle_counter_i_counter_upd_2, cs_registers_i_mcycle_counter_i_counter_upd_1, cs_registers_i_minstret_counter_i_counter_upd_63, cs_registers_i_minstret_counter_i_counter_upd_62, cs_registers_i_minstret_counter_i_counter_upd_61, cs_registers_i_minstret_counter_i_counter_upd_60, cs_registers_i_minstret_counter_i_counter_upd_59, cs_registers_i_minstret_counter_i_counter_upd_58, cs_registers_i_minstret_counter_i_counter_upd_57, cs_registers_i_minstret_counter_i_counter_upd_56, cs_registers_i_minstret_counter_i_counter_upd_55, cs_registers_i_minstret_counter_i_counter_upd_54, cs_registers_i_minstret_counter_i_counter_upd_53, cs_registers_i_minstret_counter_i_counter_upd_52, cs_registers_i_minstret_counter_i_counter_upd_51, cs_registers_i_minstret_counter_i_counter_upd_50, cs_registers_i_minstret_counter_i_counter_upd_49, cs_registers_i_minstret_counter_i_counter_upd_48, cs_registers_i_minstret_counter_i_counter_upd_47, cs_registers_i_minstret_counter_i_counter_upd_46, cs_registers_i_minstret_counter_i_counter_upd_45, cs_registers_i_minstret_counter_i_counter_upd_44, cs_registers_i_minstret_counter_i_counter_upd_43, cs_registers_i_minstret_counter_i_counter_upd_42, cs_registers_i_minstret_counter_i_counter_upd_41, cs_registers_i_minstret_counter_i_counter_upd_40, cs_registers_i_minstret_counter_i_counter_upd_39, cs_registers_i_minstret_counter_i_counter_upd_38, cs_registers_i_minstret_counter_i_counter_upd_37, cs_registers_i_minstret_counter_i_counter_upd_36, cs_registers_i_minstret_counter_i_counter_upd_35, cs_registers_i_minstret_counter_i_counter_upd_34, cs_registers_i_minstret_counter_i_counter_upd_33, cs_registers_i_minstret_counter_i_counter_upd_32, cs_registers_i_minstret_counter_i_counter_upd_31, cs_registers_i_minstret_counter_i_counter_upd_30, cs_registers_i_minstret_counter_i_counter_upd_29, cs_registers_i_minstret_counter_i_counter_upd_28, cs_registers_i_minstret_counter_i_counter_upd_27, cs_registers_i_minstret_counter_i_counter_upd_26, cs_registers_i_minstret_counter_i_counter_upd_25, cs_registers_i_minstret_counter_i_counter_upd_24, cs_registers_i_minstret_counter_i_counter_upd_23, cs_registers_i_minstret_counter_i_counter_upd_22, cs_registers_i_minstret_counter_i_counter_upd_21, cs_registers_i_minstret_counter_i_counter_upd_20, cs_registers_i_minstret_counter_i_counter_upd_19, cs_registers_i_minstret_counter_i_counter_upd_18, cs_registers_i_minstret_counter_i_counter_upd_17, cs_registers_i_minstret_counter_i_counter_upd_16, cs_registers_i_minstret_counter_i_counter_upd_15, cs_registers_i_minstret_counter_i_counter_upd_14, cs_registers_i_minstret_counter_i_counter_upd_13, cs_registers_i_minstret_counter_i_counter_upd_12, cs_registers_i_minstret_counter_i_counter_upd_11, cs_registers_i_minstret_counter_i_counter_upd_10, cs_registers_i_minstret_counter_i_counter_upd_9, cs_registers_i_minstret_counter_i_counter_upd_8, cs_registers_i_minstret_counter_i_counter_upd_7, cs_registers_i_minstret_counter_i_counter_upd_6, cs_registers_i_minstret_counter_i_counter_upd_5, cs_registers_i_minstret_counter_i_counter_upd_4, cs_registers_i_minstret_counter_i_counter_upd_3, cs_registers_i_minstret_counter_i_counter_upd_2, cs_registers_i_minstret_counter_i_counter_upd_1, n16336, n19748, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n10550, n10552, n10554, n10556, n10558, n10560, n10562, n10564, n10566, n10568, n10570, n10572, n10574, n10576, n10578, n10580, n10582, n10584, n10586, n10588, n10590, n10592, n10594, n10596, n10598, n10600, n10602, n10604, n10606, n10608, n10610, n10612, n10613, n10615, n10617, n10621, n10622, n10623, n10625, n10626, n10627, n10628, n10629, n10631, n10632, n10633, n10635, n10636, n10637, n10644, n15928, n10646, n10647, n10648, n10650, n10651, n10652, n10653, n10654, n10655, n10661, n10662, n10663, n10665, n10666, n10667, n10669, n10670, n10671, n10673, n10674, n10675, n10677, n10679, n10680, n10681, n10683, n10684, n10685, n10686, n10692, n10693, n10694, n10695, n10696, n10698, n10704, n10705, n10706, n10707, n10708, n10709, n10711, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10725, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10739, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10753, n10759, n10760, n10761, n10762, n10763, n10764, n10766, n10768, n10769, n10770, n10772, n10773, n10774, n10775, n10776, n15817, n10782, n10783, n10784, n10785, n10787, n10788, n10789, n10790, n10797, n10798, n10799, n10800, n10802, n10803, n10804, n10805, n10811, n10812, n10813, n10814, n10816, n10817, n10818, n10819, n10820, n10826, n10827, n10828, n10829, n10831, n10832, n10833, n10839, n10841, n10842, n10843, n10844, n10846, n10847, n10848, n10849, n10855, n10856, n10858, n10859, n10860, n10861, n10863, n10864, n10865, n10866, n10871, n10873, n10874, n10875, n10876, n10878, n10879, n10880, n10886, n10888, n10889, n10890, n10891, n10893, n10894, n10895, n10896, n10901, n10903, n10904, n10905, n10906, n10908, n10909, n10910, n10911, n10916, n10918, n10919, n10920, n10921, n10923, n10924, n10925, n10926, n10931, n10933, n10934, n10935, n10936, n10938, n10939, n10940, n10946, n10948, n10949, n10950, n10951, n10953, n10954, n10955, n10956, n10961, n10963, n10964, n10965, n10966, n10968, n10969, n10970, n10976, n10979, n10981, n11008, n15919, n11515, n11019, n11020, n11021, n11022, n11031, n11032, n11033, n11034, n11036, n11037, n11038, n11039, n11040, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11492, n11059, n11060, n11061, n11062, n11064, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11090, n11091, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11144, n11145, n11146, n11147, n11148, n11500, n11153, n11154, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11217, n11185, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11215, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11216, n11218, n11220, n11221, n11222, n11231, n11242, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11289, n11257, n11258, n11259, n11262, n11263, n11264, n11265, n11266, n11267, n11274, n11277, n11278, n11279, n11281, n11282, n11285, n11286, n11287, n11290, n11291, n11292, n11293, n11294, n11295, n11297, n11296, n11298, n11299, n11300, n11516, n11301, n11498, n11514, n11302, n11519, n15913, n11307, n11308, n11517, n15826, n16082, n11311, n11312, n11313, n15885, n11493, n11316, n11317, n11318, n11319, n11320, n11321, n11501, n11322, n11504, n15890, n15889, n11323, n11324, n11325, n11326, n11502, n11327, n11503, n11328, n11329, n15809, n15806, n11330, n11331, n11332, n11333, n11334, n11336, n11338, n11339, n11340, n16123, n15828, n11345, n11375, n11380, n11383, n11388, n11389, n11391, n11392, n11394, n11396, n11397, n11399, n11400, n11406, n11458, n11459, n11460, n11464, n11465, n11466, n11467, n11469, n11471, n11475, n11478, n11509, n11479, n11480, n11482, n11483, n11485, n11488, n11489, n11490, n11491, n11495, n11496, n11499, n11505, n11506, n11508, n11510, n11512, n11513;
NAND2_X4 U5641 ( .A1(n5584), .A2(n5585), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9) );
NAND2_X4 U5644 ( .A1(n5587), .A2(n5588), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8) );
NAND2_X4 U5647 ( .A1(n5589), .A2(n5590), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7) );
NAND2_X4 U5650 ( .A1(n5591), .A2(n5592), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6) );
NAND2_X4 U5653 ( .A1(n5593), .A2(n5594), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5) );
NAND2_X4 U5656 ( .A1(n5595), .A2(n5596), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4) );
NAND2_X4 U5659 ( .A1(n5597), .A2(n5598), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3) );
NAND2_X4 U5662 ( .A1(n5599), .A2(n5600), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2) );
NAND2_X4 U5665 ( .A1(n5601), .A2(n5602), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1) );
NAND2_X4 U5668 ( .A1(n5603), .A2(n5604), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15) );
NAND2_X4 U5677 ( .A1(n5609), .A2(n5610), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12) );
NAND2_X4 U5680 ( .A1(n5611), .A2(n5612), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11) );
NAND2_X4 U5683 ( .A1(n5613), .A2(n5614), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10) );
NAND2_X4 U5712 ( .A1(n5631), .A2(n5632), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2) );
NOR2_X2 U15105 ( .A1(n6222), .A2(n20961), .ZN(n5916) ); 
NAND2_X1 U15106 ( .A1(n6227), .A2(n6222), .ZN(n5917) );
NOR2_X1 U15107 ( .A1(n33), .A2(n1049), .ZN(n49) );
NOR2_X2 U15108 ( .A1(n2058), .A2(n16454), .ZN(n2142) );
INV_X4 U15109 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_1), .ZN(n20675) );
NAND2_X2 U15110 ( .A1(n5633), .A2(n5634), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_1) );
INV_X2 U15111 ( .A(n23144), .ZN(n20620) );
OR2_X1 U15112 ( .A1(n1317), .A2(n1318), .ZN(n15794) );
AND2_X1 U15113 ( .A1(n1315), .A2(n20819), .ZN(n15795) );
AND2_X1 U15114 ( .A1(n9923), .A2(n20825), .ZN(n15796) );
AND2_X1 U15115 ( .A1(alu_adder_result_ex_0), .A2(alu_adder_result_ex_1), .ZN(n15797) );
OR2_X1 U15116 ( .A1(n1318), .A2(n1319), .ZN(n15801) );
AND2_X1 U15117 ( .A1(alu_adder_result_ex_1), .A2(n20757), .ZN(n15802) );
AND2_X1 U15118 ( .A1(n7569), .A2(n7570), .ZN(n15808) );
OR2_X1 U15119 ( .A1(n4958), .A2(n20921), .ZN(n15811) );
AND2_X1 U15120 ( .A1(n5777), .A2(n5778), .ZN(n15829) );
AND2_X1 U15121 ( .A1(n5773), .A2(n5774), .ZN(n15830) );
AND2_X1 U15122 ( .A1(n5779), .A2(n5780), .ZN(n15831) );
AND2_X1 U15123 ( .A1(n5791), .A2(n5792), .ZN(n15832) );
AND2_X1 U15124 ( .A1(n5767), .A2(n5768), .ZN(n15833) );
AND2_X1 U15125 ( .A1(n5759), .A2(n5760), .ZN(n15834) );
AND2_X1 U15126 ( .A1(n5751), .A2(n5752), .ZN(n15835) );
AND2_X1 U15127 ( .A1(n5769), .A2(n5770), .ZN(n15836) );
AND2_X1 U15128 ( .A1(n5761), .A2(n5762), .ZN(n15837) );
AND2_X1 U15129 ( .A1(n5755), .A2(n5756), .ZN(n15838) );
AND2_X1 U15130 ( .A1(n5771), .A2(n5772), .ZN(n15839) );
AND2_X1 U15131 ( .A1(n5763), .A2(n5764), .ZN(n15840) );
AND2_X1 U15132 ( .A1(n5757), .A2(n5758), .ZN(n15841) );
AND2_X1 U15133 ( .A1(n5765), .A2(n5766), .ZN(n15842) );
AND2_X1 U15134 ( .A1(n5743), .A2(n5744), .ZN(n15843) );
AND2_X1 U15135 ( .A1(n5745), .A2(n5746), .ZN(n15844) );
AND2_X1 U15136 ( .A1(n5747), .A2(n5748), .ZN(n15845) );
AND2_X1 U15137 ( .A1(n5749), .A2(n5750), .ZN(n15846) );
AND2_X1 U15138 ( .A1(n5785), .A2(n5786), .ZN(n15847) );
AND2_X1 U15139 ( .A1(n5793), .A2(n5794), .ZN(n15848) );
AND2_X1 U15140 ( .A1(n5787), .A2(n5788), .ZN(n15849) );
AND2_X1 U15141 ( .A1(n5789), .A2(n5790), .ZN(n15850) );
AND2_X1 U15142 ( .A1(n5781), .A2(n5782), .ZN(n15851) );
AND2_X1 U15143 ( .A1(n5783), .A2(n5784), .ZN(n15852) );
AND2_X1 U15144 ( .A1(n5741), .A2(n5742), .ZN(n15853) );
AND2_X1 U15145 ( .A1(n5795), .A2(n5796), .ZN(n15854) );
AND2_X1 U15146 ( .A1(n5737), .A2(n5738), .ZN(n15855) );
AND2_X1 U15147 ( .A1(n5739), .A2(n5740), .ZN(n15856) );
AND2_X1 U15148 ( .A1(n21999), .A2(n21998), .ZN(n15857) );
NAND2_X1 U15149 ( .A1(n20855), .A2(n20850), .ZN(n22074) );
NAND2_X1 U15150 ( .A1(n20863), .A2(n20856), .ZN(n21946) );
BUF_X1 U15151 ( .A(n4067), .Z(n16425) );
NOR2_X1 U15152 ( .A1(n21231), .A2(n21230), .ZN(alu_adder_result_ex_1) );
INV_X1 U15153 ( .A(ex_block_i_alu_i_shift_amt_4), .ZN(n20850) );
NAND2_X1 U15154 ( .A1(ex_block_i_alu_i_shift_amt_4), .A2(ex_block_i_alu_i_N294), .ZN(n21999) );
OR2_X1 U15155 ( .A1(n21960), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n22078) );
NOR2_X1 U15156 ( .A1(n6303), .A2(n6304), .ZN(ex_block_i_alu_i_N294) );
NAND2_X1 U15157 ( .A1(ex_block_i_alu_i_shift_amt_2), .A2(n20856), .ZN(n21960) );
BUF_X1 U15158 ( .A(n5386), .Z(n16413) );
INV_X1 U15159 ( .A(n16262), .ZN(n16391) );
INV_X1 U15160 ( .A(n16262), .ZN(n16390) );
INV_X1 U15161 ( .A(alu_operand_b_ex_4), .ZN(n20853) );
NOR2_X1 U15162 ( .A1(n20871), .A2(alu_operand_b_ex_1), .ZN(n7571) );
NOR2_X1 U15163 ( .A1(n5120), .A2(n5127), .ZN(n7581) );
BUF_X1 U15164 ( .A(n1708), .Z(n16458) );
NAND2_X1 U15165 ( .A1(n5800), .A2(n5801), .ZN(ex_block_i_alu_i_shift_amt_4) );
NAND2_X1 U15166 ( .A1(n1365), .A2(n1366), .ZN(n16335) );
NOR2_X1 U15167 ( .A1(n2727), .A2(n19942), .ZN(n2112) );
NOR2_X1 U15168 ( .A1(n5090), .A2(n1431), .ZN(n4417) );
NOR2_X1 U15169 ( .A1(n15818), .A2(n16115), .ZN(n1039) );
NOR2_X1 U15170 ( .A1(n2727), .A2(n2432), .ZN(n2270) );
NAND2_X1 U15171 ( .A1(n10494), .A2(n10495), .ZN(alu_operand_b_ex_1) );
NAND2_X1 U15172 ( .A1(n10028), .A2(n10029), .ZN(n1297) );
AND2_X1 U15173 ( .A1(n19967), .A2(n1048), .ZN(n367) );
NAND2_X1 U15174 ( .A1(n11460), .A2(crash_dump_o_65_), .ZN(n2782) );
NOR2_X1 U15175 ( .A1(n1058), .A2(n11064), .ZN(n163) );
NAND2_X1 U15176 ( .A1(n5710), .A2(n20992), .ZN(n5687) );
NOR2_X1 U15177 ( .A1(n3721), .A2(n11475), .ZN(n3019) );
NAND2_X1 U15178 ( .A1(n10448), .A2(n11520), .ZN(n1431) );
NAND2_X1 U15179 ( .A1(n2844), .A2(n2845), .ZN(n2042) );
NOR2_X1 U15180 ( .A1(instr_err_i), .A2(n15920), .ZN(n2753) );
NAND2_X1 U15181 ( .A1(n11500), .A2(n15907), .ZN(n1444) );
INV_X1 U15182 ( .A(n23496), .ZN(n16198) );
INV_X1 U15183 ( .A(n23635), .ZN(n16199) );
INV_X2 U15184 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n16200) );
INV_X1 U15185 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n20683) );
BUF_X1 U15186 ( .A(n19883), .Z(n16345) );
INV_X1 U15187 ( .A(n15801), .ZN(n16474) );
INV_X1 U15188 ( .A(n15801), .ZN(n16475) );
INV_X1 U15189 ( .A(n15795), .ZN(n16473) );
INV_X1 U15190 ( .A(n15794), .ZN(n16472) );
INV_X1 U15191 ( .A(n16455), .ZN(n16451) );
INV_X1 U15192 ( .A(n16456), .ZN(n16452) );
INV_X1 U15193 ( .A(n16457), .ZN(n16453) );
INV_X1 U15194 ( .A(n16456), .ZN(n16450) );
INV_X1 U15195 ( .A(n3054), .ZN(n19883) );
INV_X1 U15196 ( .A(ex_block_i_alu_is_equal_result), .ZN(n20111) );
NOR2_X1 U15197 ( .A1(n20172), .A2(n20926), .ZN(n3747) );
NOR2_X1 U15198 ( .A1(n20404), .A2(n20926), .ZN(n3820) );
NOR2_X1 U15199 ( .A1(n20326), .A2(n20926), .ZN(n3797) );
NOR2_X1 U15200 ( .A1(n20210), .A2(n20926), .ZN(n3758) );
NOR2_X1 U15201 ( .A1(n16469), .A2(n20365), .ZN(n677) );
NOR2_X1 U15202 ( .A1(n16469), .A2(n20326), .ZN(n639) );
NOR2_X1 U15203 ( .A1(n16469), .A2(n20287), .ZN(n599) );
NOR2_X1 U15204 ( .A1(n90), .A2(n20248), .ZN(n559) );
NOR2_X1 U15205 ( .A1(n90), .A2(n20210), .ZN(n519) );
NOR2_X1 U15206 ( .A1(n90), .A2(n20172), .ZN(n436) );
NOR2_X1 U15207 ( .A1(n20641), .A2(n20926), .ZN(n3887) );
NOR2_X1 U15208 ( .A1(n20603), .A2(n20926), .ZN(n3876) );
NOR2_X1 U15209 ( .A1(n20523), .A2(n20926), .ZN(n3853) );
NOR2_X1 U15210 ( .A1(n20483), .A2(n20926), .ZN(n3842) );
NOR2_X1 U15211 ( .A1(n20443), .A2(n20926), .ZN(n3831) );
NOR2_X1 U15212 ( .A1(n90), .A2(n20603), .ZN(n948) );
NOR2_X1 U15213 ( .A1(n90), .A2(n20563), .ZN(n867) );
NOR2_X1 U15214 ( .A1(n90), .A2(n20523), .ZN(n828) );
NOR2_X1 U15215 ( .A1(n90), .A2(n20483), .ZN(n790) );
NOR2_X1 U15216 ( .A1(n90), .A2(n20443), .ZN(n752) );
NOR2_X1 U15217 ( .A1(n90), .A2(n20404), .ZN(n715) );
NOR2_X1 U15218 ( .A1(n20696), .A2(n20926), .ZN(n3943) );
NOR2_X1 U15219 ( .A1(n20692), .A2(n20926), .ZN(n3932) );
NOR2_X1 U15220 ( .A1(n20688), .A2(n20926), .ZN(n3921) );
NOR2_X1 U15221 ( .A1(n20676), .A2(n20926), .ZN(n3898) );
NOR2_X1 U15222 ( .A1(n90), .A2(n20684), .ZN(n1084) );
NOR2_X1 U15223 ( .A1(n90), .A2(n20676), .ZN(n1025) );
NOR2_X1 U15224 ( .A1(n90), .A2(n20641), .ZN(n987) );
INV_X1 U15225 ( .A(n87), .ZN(n20818) );
BUF_X1 U15226 ( .A(n90), .Z(n16469) );
BUF_X1 U15227 ( .A(n15801), .Z(n16476) );
BUF_X1 U15228 ( .A(n83), .Z(n16470) );
INV_X1 U15229 ( .A(n15796), .ZN(n16361) );
BUF_X1 U15230 ( .A(n1566), .Z(n16462) );
INV_X1 U15231 ( .A(n16363), .ZN(n16362) );
INV_X1 U15232 ( .A(n15797), .ZN(n16463) );
INV_X1 U15233 ( .A(n15802), .ZN(n16407) );
INV_X1 U15234 ( .A(n15797), .ZN(n16464) );
INV_X1 U15235 ( .A(n15802), .ZN(n16406) );
INV_X1 U15236 ( .A(n8118), .ZN(n20859) );
BUF_X1 U15237 ( .A(n8437), .Z(n16378) );
BUF_X1 U15238 ( .A(n8150), .Z(n16381) );
BUF_X1 U15239 ( .A(n7318), .Z(n16396) );
BUF_X1 U15240 ( .A(n8169), .Z(n16380) );
BUF_X1 U15241 ( .A(n19977), .Z(n16349) );
BUF_X1 U15242 ( .A(n19977), .Z(n16348) );
BUF_X1 U15243 ( .A(n3396), .Z(n16432) );
BUF_X1 U15244 ( .A(n19976), .Z(n16347) );
NAND2_X1 U15245 ( .A1(n16440), .A2(n16456), .ZN(n3054) );
BUF_X1 U15246 ( .A(n6552), .Z(n16404) );
BUF_X1 U15247 ( .A(n16457), .Z(n16455) );
BUF_X1 U15248 ( .A(n16457), .Z(n16456) );
BUF_X1 U15249 ( .A(n16457), .Z(n16454) );
NOR2_X1 U15250 ( .A1(n21648), .A2(n21647), .ZN(ex_block_i_alu_is_equal_result) );
NAND2_X1 U15251 ( .A1(n21646), .A2(n21645), .ZN(n21647) );
NOR2_X1 U15252 ( .A1(n21638), .A2(n21637), .ZN(n21646) );
INV_X1 U15253 ( .A(data_addr_o_30_), .ZN(n20172) );
NOR2_X1 U15254 ( .A1(n20112), .A2(n20926), .ZN(n3734) );
NOR2_X1 U15255 ( .A1(data_addr_o_27_), .A2(data_addr_o_26_), .ZN(n21621) );
NOR2_X1 U15256 ( .A1(data_addr_o_29_), .A2(data_addr_o_28_), .ZN(n21620) );
NOR2_X1 U15257 ( .A1(n16469), .A2(n20112), .ZN(n391) );
NOR2_X1 U15258 ( .A1(n21624), .A2(n21623), .ZN(n21632) );
NAND2_X1 U15259 ( .A1(n21622), .A2(n21621), .ZN(n21623) );
NAND2_X1 U15260 ( .A1(n21620), .A2(n21619), .ZN(n21624) );
NOR2_X1 U15261 ( .A1(data_addr_o_25_), .A2(data_addr_o_24_), .ZN(n21622) );
INV_X1 U15262 ( .A(data_addr_o_26_), .ZN(n20326) );
INV_X1 U15263 ( .A(data_addr_o_24_), .ZN(n20404) );
INV_X1 U15264 ( .A(data_addr_o_29_), .ZN(n20210) );
INV_X1 U15265 ( .A(data_addr_o_27_), .ZN(n20287) );
INV_X1 U15266 ( .A(data_addr_o_25_), .ZN(n20365) );
INV_X1 U15267 ( .A(data_addr_o_28_), .ZN(n20248) );
NOR2_X1 U15268 ( .A1(data_addr_o_23_), .A2(data_addr_o_22_), .ZN(n21639) );
NOR2_X1 U15269 ( .A1(n21644), .A2(n21643), .ZN(n21645) );
NAND2_X1 U15270 ( .A1(n21642), .A2(n21641), .ZN(n21643) );
NAND2_X1 U15271 ( .A1(n21640), .A2(n21639), .ZN(n21644) );
NOR2_X1 U15272 ( .A1(data_addr_o_18_), .A2(data_addr_o_17_), .ZN(n21642) );
NOR2_X1 U15273 ( .A1(data_addr_o_21_), .A2(data_addr_o_20_), .ZN(n21640) );
INV_X1 U15274 ( .A(data_addr_o_22_), .ZN(n20483) );
INV_X1 U15275 ( .A(data_addr_o_19_), .ZN(n20603) );
INV_X1 U15276 ( .A(data_addr_o_23_), .ZN(n20443) );
INV_X1 U15277 ( .A(data_addr_o_21_), .ZN(n20523) );
INV_X1 U15278 ( .A(data_addr_o_18_), .ZN(n20641) );
INV_X1 U15279 ( .A(data_addr_o_20_), .ZN(n20563) );
NAND2_X1 U15280 ( .A1(n21634), .A2(n21633), .ZN(n21638) );
NOR2_X1 U15281 ( .A1(data_addr_o_14_), .A2(data_addr_o_13_), .ZN(n21634) );
NOR2_X1 U15282 ( .A1(data_addr_o_16_), .A2(data_addr_o_15_), .ZN(n21633) );
INV_X1 U15283 ( .A(data_addr_o_17_), .ZN(n20676) );
INV_X1 U15284 ( .A(data_addr_o_15_), .ZN(n20688) );
INV_X1 U15285 ( .A(data_addr_o_13_), .ZN(n20696) );
INV_X1 U15286 ( .A(data_addr_o_14_), .ZN(n20692) );
NOR2_X1 U15287 ( .A1(n20700), .A2(n20926), .ZN(n3954) );
INV_X1 U15288 ( .A(data_addr_o_16_), .ZN(n20684) );
NOR2_X2 U15289 ( .A1(n16466), .A2(n1318), .ZN(n87) );
INV_X1 U15290 ( .A(n1334), .ZN(n20821) );
INV_X1 U15291 ( .A(n3018), .ZN(n16439) );
NOR2_X1 U15292 ( .A1(n20818), .A2(n16247), .ZN(n394) );
NOR2_X1 U15293 ( .A1(n20727), .A2(n20926), .ZN(n4021) );
NOR2_X1 U15294 ( .A1(n20721), .A2(n20926), .ZN(n4013) );
NOR2_X1 U15295 ( .A1(n20716), .A2(n20926), .ZN(n3999) );
NOR2_X1 U15296 ( .A1(n20708), .A2(n20926), .ZN(n3977) );
NOR2_X1 U15297 ( .A1(n20712), .A2(n20926), .ZN(n3988) );
INV_X1 U15298 ( .A(n8624), .ZN(n16363) );
INV_X1 U15299 ( .A(n1318), .ZN(n20819) );
NAND2_X1 U15300 ( .A1(n1342), .A2(n20819), .ZN(n90) );
NAND2_X1 U15301 ( .A1(n9982), .A2(n9983), .ZN(n9981) );
NOR2_X1 U15302 ( .A1(n16384), .A2(n16363), .ZN(n9983) );
NOR2_X1 U15303 ( .A1(n16386), .A2(n16201), .ZN(n9982) );
INV_X1 U15304 ( .A(n16201), .ZN(n16367) );
INV_X1 U15305 ( .A(n16201), .ZN(n16368) );
BUF_X1 U15306 ( .A(n8590), .Z(n16370) );
BUF_X1 U15307 ( .A(n8591), .Z(n16369) );
BUF_X1 U15308 ( .A(n20866), .Z(n16351) );
NAND2_X1 U15309 ( .A1(n16361), .A2(n8575), .ZN(n8758) );
BUF_X1 U15310 ( .A(n6318), .Z(n16405) );
BUF_X1 U15311 ( .A(n8585), .Z(n16371) );
BUF_X1 U15312 ( .A(n8576), .Z(n16373) );
INV_X1 U15313 ( .A(n16384), .ZN(n16383) );
INV_X1 U15314 ( .A(n21946), .ZN(n20855) );
INV_X1 U15315 ( .A(n22074), .ZN(n20849) );
NAND2_X1 U15316 ( .A1(n20868), .A2(n20860), .ZN(n8118) );
NAND2_X1 U15317 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_30), .A2(n87), .ZN(n908) );
NAND2_X1 U15318 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_29), .A2(n87), .ZN(n477) );
NAND2_X1 U15319 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_28), .A2(n87), .ZN(n347) );
NAND2_X1 U15320 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_27), .A2(n87), .ZN(n306) );
NOR2_X1 U15321 ( .A1(n20642), .A2(n22074), .ZN(n21867) );
NOR2_X1 U15322 ( .A1(n20677), .A2(n22074), .ZN(n21858) );
NOR2_X1 U15323 ( .A1(n20643), .A2(n22074), .ZN(n21832) );
NOR2_X1 U15324 ( .A1(n20605), .A2(n22074), .ZN(n21813) );
NOR2_X1 U15325 ( .A1(n20565), .A2(n22074), .ZN(n21786) );
NOR2_X1 U15326 ( .A1(n20525), .A2(n22074), .ZN(n21744) );
NOR2_X1 U15327 ( .A1(n20484), .A2(n22074), .ZN(n22077) );
NOR2_X1 U15328 ( .A1(n20444), .A2(n22074), .ZN(n22067) );
NOR2_X1 U15329 ( .A1(n20749), .A2(n20926), .ZN(n3727) );
NOR2_X1 U15330 ( .A1(n20743), .A2(n20926), .ZN(n4045) );
NOR2_X1 U15331 ( .A1(n20738), .A2(n20926), .ZN(n4037) );
NOR2_X1 U15332 ( .A1(n20732), .A2(n20926), .ZN(n4029) );
NOR2_X1 U15333 ( .A1(n16470), .A2(n20127), .ZN(n1076) );
INV_X1 U15334 ( .A(ex_block_i_alu_i_shift_result_ext_signed_16), .ZN(n20127) );
NOR2_X1 U15335 ( .A1(n20604), .A2(n21946), .ZN(n21680) );
NOR2_X1 U15336 ( .A1(n20327), .A2(n21946), .ZN(n21947) );
NOR2_X1 U15337 ( .A1(n20366), .A2(n21946), .ZN(n21940) );
NOR2_X1 U15338 ( .A1(n20405), .A2(n21946), .ZN(n21934) );
NOR2_X1 U15339 ( .A1(n20445), .A2(n21946), .ZN(n21927) );
NOR2_X1 U15340 ( .A1(n20485), .A2(n21946), .ZN(n21892) );
NOR2_X1 U15341 ( .A1(n20524), .A2(n21946), .ZN(n21883) );
NOR2_X1 U15342 ( .A1(n20564), .A2(n21946), .ZN(n21874) );
NOR2_X1 U15343 ( .A1(n83), .A2(n20126), .ZN(n1018) );
INV_X1 U15344 ( .A(ex_block_i_alu_i_shift_result_ext_signed_17), .ZN(n20126) );
NOR2_X1 U15345 ( .A1(n83), .A2(n20125), .ZN(n980) );
INV_X1 U15346 ( .A(ex_block_i_alu_i_shift_result_ext_signed_18), .ZN(n20125) );
NOR2_X1 U15347 ( .A1(n83), .A2(n20124), .ZN(n941) );
INV_X1 U15348 ( .A(ex_block_i_alu_i_shift_result_ext_signed_19), .ZN(n20124) );
NOR2_X1 U15349 ( .A1(n83), .A2(n20123), .ZN(n860) );
INV_X1 U15350 ( .A(ex_block_i_alu_i_shift_result_ext_signed_20), .ZN(n20123) );
NOR2_X1 U15351 ( .A1(n83), .A2(n20122), .ZN(n821) );
INV_X1 U15352 ( .A(ex_block_i_alu_i_shift_result_ext_signed_21), .ZN(n20122) );
NOR2_X1 U15353 ( .A1(n83), .A2(n20120), .ZN(n745) );
INV_X1 U15354 ( .A(ex_block_i_alu_i_shift_result_ext_signed_23), .ZN(n20120) );
NOR2_X1 U15355 ( .A1(n83), .A2(n20119), .ZN(n708) );
INV_X1 U15356 ( .A(ex_block_i_alu_i_shift_result_ext_signed_24), .ZN(n20119) );
NOR2_X1 U15357 ( .A1(n83), .A2(n20118), .ZN(n670) );
INV_X1 U15358 ( .A(ex_block_i_alu_i_shift_result_ext_signed_25), .ZN(n20118) );
NOR2_X1 U15359 ( .A1(n83), .A2(n20117), .ZN(n631) );
INV_X1 U15360 ( .A(ex_block_i_alu_i_shift_result_ext_signed_26), .ZN(n20117) );
NOR2_X1 U15361 ( .A1(n83), .A2(n20116), .ZN(n591) );
INV_X1 U15362 ( .A(ex_block_i_alu_i_shift_result_ext_signed_27), .ZN(n20116) );
NOR2_X1 U15363 ( .A1(n16470), .A2(n20115), .ZN(n551) );
INV_X1 U15364 ( .A(ex_block_i_alu_i_shift_result_ext_signed_28), .ZN(n20115) );
NOR2_X1 U15365 ( .A1(n16470), .A2(n20114), .ZN(n511) );
INV_X1 U15366 ( .A(ex_block_i_alu_i_shift_result_ext_signed_29), .ZN(n20114) );
NOR2_X1 U15367 ( .A1(n16470), .A2(n20113), .ZN(n428) );
INV_X1 U15368 ( .A(ex_block_i_alu_i_shift_result_ext_signed_30), .ZN(n20113) );
NOR2_X1 U15369 ( .A1(n20121), .A2(n16470), .ZN(n783) );
INV_X1 U15370 ( .A(ex_block_i_alu_i_shift_result_ext_signed_22), .ZN(n20121) );
INV_X1 U15371 ( .A(n21810), .ZN(n20133) );
INV_X1 U15372 ( .A(n21876), .ZN(n20131) );
NAND2_X1 U15373 ( .A1(n20753), .A2(n20757), .ZN(n1566) );
INV_X1 U15374 ( .A(n9868), .ZN(n20843) );
INV_X1 U15375 ( .A(n9907), .ZN(n20823) );
OR2_X1 U15376 ( .A1(n1335), .A2(n1318), .ZN(n83) );
INV_X1 U15377 ( .A(n6561), .ZN(n19971) );
INV_X1 U15378 ( .A(n7257), .ZN(n19973) );
INV_X1 U15379 ( .A(n16442), .ZN(n16440) );
BUF_X1 U15380 ( .A(n20909), .Z(n16352) );
INV_X1 U15381 ( .A(n15808), .ZN(n16394) );
INV_X1 U15382 ( .A(n15808), .ZN(n16393) );
BUF_X1 U15383 ( .A(n4061), .Z(n16427) );
BUF_X1 U15384 ( .A(n7178), .Z(n16397) );
BUF_X1 U15385 ( .A(n7178), .Z(n16398) );
INV_X1 U15386 ( .A(n16442), .ZN(n16441) );
BUF_X1 U15387 ( .A(n8149), .Z(n16382) );
INV_X1 U15388 ( .A(n2117), .ZN(n19875) );
NOR2_X1 U15389 ( .A1(n6698), .A2(n8118), .ZN(n7078) );
INV_X1 U15390 ( .A(n3611), .ZN(n16430) );
NOR2_X1 U15391 ( .A1(n7562), .A2(n15808), .ZN(n7318) );
NOR2_X1 U15392 ( .A1(n16442), .A2(n19883), .ZN(n3396) );
NAND2_X1 U15393 ( .A1(n6561), .A2(n16404), .ZN(n6554) );
INV_X1 U15394 ( .A(n8883), .ZN(n19982) );
INV_X1 U15395 ( .A(n2036), .ZN(n19878) );
NOR2_X1 U15396 ( .A1(n19805), .A2(n16378), .ZN(n8643) );
NOR2_X1 U15397 ( .A1(n20712), .A2(n4067), .ZN(n4063) );
NOR2_X1 U15398 ( .A1(n20716), .A2(n4067), .ZN(n4071) );
NOR2_X1 U15399 ( .A1(n20721), .A2(n4067), .ZN(n4077) );
NOR2_X1 U15400 ( .A1(n20727), .A2(n4067), .ZN(n4083) );
NOR2_X1 U15401 ( .A1(n20732), .A2(n4067), .ZN(n4089) );
NOR2_X1 U15402 ( .A1(n20738), .A2(n4067), .ZN(n4095) );
NOR2_X1 U15403 ( .A1(n20743), .A2(n4067), .ZN(n4101) );
NOR2_X1 U15404 ( .A1(n20112), .A2(n4067), .ZN(n4107) );
NOR2_X1 U15405 ( .A1(n19803), .A2(n16381), .ZN(n8228) );
NOR2_X1 U15406 ( .A1(n19803), .A2(n16378), .ZN(n8515) );
NOR2_X1 U15407 ( .A1(n19805), .A2(n16381), .ZN(n8272) );
NOR2_X1 U15408 ( .A1(n20753), .A2(n4067), .ZN(n4185) );
INV_X1 U15409 ( .A(n16429), .ZN(n16431) );
NOR2_X1 U15410 ( .A1(n19809), .A2(n8150), .ZN(n8368) );
NOR2_X1 U15411 ( .A1(n19809), .A2(n8437), .ZN(n9385) );
NOR2_X1 U15412 ( .A1(n20172), .A2(n16425), .ZN(n4113) );
NOR2_X1 U15413 ( .A1(n20749), .A2(n16425), .ZN(n4119) );
NOR2_X1 U15414 ( .A1(n20210), .A2(n16425), .ZN(n4125) );
NOR2_X1 U15415 ( .A1(n20248), .A2(n16425), .ZN(n4131) );
NOR2_X1 U15416 ( .A1(n20287), .A2(n16425), .ZN(n4137) );
NOR2_X1 U15417 ( .A1(n20326), .A2(n16425), .ZN(n4143) );
NOR2_X1 U15418 ( .A1(n20365), .A2(n16425), .ZN(n4149) );
NOR2_X1 U15419 ( .A1(n20404), .A2(n16425), .ZN(n4155) );
NOR2_X1 U15420 ( .A1(n20443), .A2(n16425), .ZN(n4161) );
NOR2_X1 U15421 ( .A1(n20483), .A2(n16425), .ZN(n4167) );
NOR2_X1 U15422 ( .A1(n20523), .A2(n16425), .ZN(n4173) );
NOR2_X1 U15423 ( .A1(n20563), .A2(n16425), .ZN(n4179) );
NOR2_X1 U15424 ( .A1(n20603), .A2(n4067), .ZN(n4191) );
NOR2_X1 U15425 ( .A1(n20641), .A2(n4067), .ZN(n4197) );
NOR2_X1 U15426 ( .A1(n20676), .A2(n4067), .ZN(n4203) );
NOR2_X1 U15427 ( .A1(n20684), .A2(n16425), .ZN(n4209) );
NOR2_X1 U15428 ( .A1(n20688), .A2(n4067), .ZN(n4215) );
NOR2_X1 U15429 ( .A1(n20692), .A2(n16425), .ZN(n4221) );
NOR2_X1 U15430 ( .A1(n20696), .A2(n4067), .ZN(n4227) );
NOR2_X1 U15431 ( .A1(n20700), .A2(n16425), .ZN(n4233) );
NOR2_X1 U15432 ( .A1(n20704), .A2(n4067), .ZN(n4239) );
NOR2_X1 U15433 ( .A1(n20708), .A2(n16425), .ZN(n4245) );
NOR2_X1 U15434 ( .A1(n20757), .A2(n4067), .ZN(n4253) );
NOR2_X1 U15435 ( .A1(n19809), .A2(n16380), .ZN(n8300) );
NOR2_X1 U15436 ( .A1(n19809), .A2(n8456), .ZN(n8877) );
NOR2_X1 U15437 ( .A1(n19803), .A2(n16380), .ZN(n8288) );
NOR2_X1 U15438 ( .A1(n19803), .A2(n8456), .ZN(n8776) );
NOR2_X1 U15439 ( .A1(n19805), .A2(n16380), .ZN(n8292) );
NOR2_X1 U15440 ( .A1(n19805), .A2(n16377), .ZN(n8822) );
NAND2_X1 U15441 ( .A1(n6190), .A2(n6186), .ZN(n10482) );
INV_X1 U15442 ( .A(n7725), .ZN(n19976) );
NOR2_X1 U15443 ( .A1(n19895), .A2(n2648), .ZN(n2647) );
OR2_X1 U15444 ( .A1(n2649), .A2(n2025), .ZN(n2648) );
NAND2_X1 U15445 ( .A1(n19979), .A2(n19980), .ZN(n8150) );
NAND2_X1 U15446 ( .A1(n19981), .A2(n19982), .ZN(n8437) );
NAND2_X1 U15447 ( .A1(n2025), .A2(n16451), .ZN(n2104) );
INV_X1 U15448 ( .A(n7803), .ZN(n19977) );
INV_X1 U15449 ( .A(n7052), .ZN(n19972) );
INV_X1 U15450 ( .A(n9891), .ZN(n19970) );
INV_X1 U15451 ( .A(n1338), .ZN(n16467) );
INV_X1 U15452 ( .A(n1338), .ZN(n16468) );
NAND2_X1 U15453 ( .A1(n2649), .A2(n16452), .ZN(n2237) );
INV_X1 U15454 ( .A(n3773), .ZN(n20926) );
INV_X1 U15455 ( .A(n3774), .ZN(n20927) );
NAND2_X1 U15456 ( .A1(n19980), .A2(n8165), .ZN(n8169) );
INV_X1 U15457 ( .A(n2696), .ZN(n19939) );
INV_X1 U15458 ( .A(n4046), .ZN(n20928) );
NAND2_X1 U15459 ( .A1(n3740), .A2(n3018), .ZN(n6552) );
INV_X1 U15460 ( .A(n2470), .ZN(n19905) );
INV_X1 U15461 ( .A(n6190), .ZN(n20955) );
INV_X1 U15462 ( .A(n10481), .ZN(n20953) );
INV_X1 U15463 ( .A(n1885), .ZN(n16457) );
AND2_X1 U15464 ( .A1(n2457), .A2(n2237), .ZN(n2461) );
NOR2_X1 U15465 ( .A1(n21216), .A2(n21215), .ZN(data_addr_o_27_) );
NOR2_X1 U15466 ( .A1(n21217), .A2(n21214), .ZN(n21216) );
AND2_X1 U15467 ( .A1(n21217), .A2(n21214), .ZN(n21215) );
NAND2_X1 U15468 ( .A1(n21213), .A2(n21212), .ZN(n21214) );
NOR2_X1 U15469 ( .A1(n21225), .A2(n21224), .ZN(data_addr_o_28_) );
NOR2_X1 U15470 ( .A1(n21232), .A2(n21223), .ZN(n21225) );
AND2_X1 U15471 ( .A1(n21232), .A2(n21223), .ZN(n21224) );
NAND2_X1 U15472 ( .A1(n21222), .A2(n21221), .ZN(n21223) );
NOR2_X1 U15473 ( .A1(n21240), .A2(n21239), .ZN(data_addr_o_29_) );
NOR2_X1 U15474 ( .A1(n21241), .A2(n21238), .ZN(n21240) );
AND2_X1 U15475 ( .A1(n21241), .A2(n21238), .ZN(n21239) );
NAND2_X1 U15476 ( .A1(n21237), .A2(n21236), .ZN(n21238) );
NOR2_X1 U15477 ( .A1(n21249), .A2(n21248), .ZN(data_addr_o_30_) );
NOR2_X1 U15478 ( .A1(n21252), .A2(n21247), .ZN(n21249) );
AND2_X1 U15479 ( .A1(n21252), .A2(n21247), .ZN(n21248) );
NAND2_X1 U15480 ( .A1(n21246), .A2(n21245), .ZN(n21247) );
INV_X1 U15481 ( .A(data_addr_o_31_), .ZN(n20112) );
NOR2_X1 U15482 ( .A1(n1407), .A2(n1408), .ZN(n1381) );
NOR2_X1 U15483 ( .A1(n16466), .A2(n15857), .ZN(n1407) );
NAND2_X1 U15484 ( .A1(alu_adder_result_ex_0), .A2(n1342), .ZN(n1410) );
NOR2_X1 U15485 ( .A1(n10107), .A2(n10108), .ZN(n10106) );
NOR2_X1 U15486 ( .A1(n10109), .A2(n10110), .ZN(n10107) );
NOR2_X1 U15487 ( .A1(n10111), .A2(n10112), .ZN(n10110) );
NOR2_X1 U15488 ( .A1(n20111), .A2(n10118), .ZN(n10109) );
NOR2_X1 U15489 ( .A1(data_addr_o_30_), .A2(data_addr_o_2_), .ZN(n21619) );
NOR2_X1 U15490 ( .A1(data_addr_o_3_), .A2(data_addr_o_31_), .ZN(n21628) );
AND2_X1 U15491 ( .A1(n10085), .A2(n10086), .ZN(n1412) );
NOR2_X1 U15492 ( .A1(n10087), .A2(n10088), .ZN(n10086) );
NOR2_X1 U15493 ( .A1(n10105), .A2(n10106), .ZN(n10085) );
NOR2_X1 U15494 ( .A1(n20111), .A2(n10089), .ZN(n10088) );
NOR2_X1 U15495 ( .A1(n21630), .A2(n21629), .ZN(n21631) );
NAND2_X1 U15496 ( .A1(n21626), .A2(n21625), .ZN(n21630) );
NAND2_X1 U15497 ( .A1(n21628), .A2(n21627), .ZN(n21629) );
NOR2_X1 U15498 ( .A1(data_addr_o_7_), .A2(data_addr_o_6_), .ZN(n21626) );
OR2_X1 U15499 ( .A1(n1411), .A2(n1412), .ZN(n1409) );
NOR2_X1 U15500 ( .A1(n21198), .A2(n21197), .ZN(data_addr_o_25_) );
NOR2_X1 U15501 ( .A1(n21199), .A2(n21196), .ZN(n21198) );
AND2_X1 U15502 ( .A1(n21199), .A2(n21196), .ZN(n21197) );
NAND2_X1 U15503 ( .A1(n21195), .A2(n21194), .ZN(n21196) );
NOR2_X1 U15504 ( .A1(n21162), .A2(n21161), .ZN(data_addr_o_21_) );
NOR2_X1 U15505 ( .A1(n21163), .A2(n21160), .ZN(n21162) );
AND2_X1 U15506 ( .A1(n21163), .A2(n21160), .ZN(n21161) );
NAND2_X1 U15507 ( .A1(n21159), .A2(n21158), .ZN(n21160) );
NOR2_X1 U15508 ( .A1(n21180), .A2(n21179), .ZN(data_addr_o_23_) );
NOR2_X1 U15509 ( .A1(n21181), .A2(n21178), .ZN(n21180) );
AND2_X1 U15510 ( .A1(n21181), .A2(n21178), .ZN(n21179) );
NAND2_X1 U15511 ( .A1(n21177), .A2(n21176), .ZN(n21178) );
NOR2_X1 U15512 ( .A1(n21171), .A2(n21170), .ZN(data_addr_o_22_) );
NOR2_X1 U15513 ( .A1(n21172), .A2(n21169), .ZN(n21171) );
AND2_X1 U15514 ( .A1(n21172), .A2(n21169), .ZN(n21170) );
NAND2_X1 U15515 ( .A1(n21168), .A2(n21167), .ZN(n21169) );
NOR2_X1 U15516 ( .A1(n21189), .A2(n21188), .ZN(data_addr_o_24_) );
NOR2_X1 U15517 ( .A1(n21190), .A2(n21187), .ZN(n21189) );
AND2_X1 U15518 ( .A1(n21190), .A2(n21187), .ZN(n21188) );
NAND2_X1 U15519 ( .A1(n21186), .A2(n21185), .ZN(n21187) );
NOR2_X1 U15520 ( .A1(n21207), .A2(n21206), .ZN(data_addr_o_26_) );
NOR2_X1 U15521 ( .A1(n21208), .A2(n21205), .ZN(n21207) );
AND2_X1 U15522 ( .A1(n21208), .A2(n21205), .ZN(n21206) );
NAND2_X1 U15523 ( .A1(n21204), .A2(n21203), .ZN(n21205) );
NOR2_X1 U15524 ( .A1(n21112), .A2(n21111), .ZN(data_addr_o_16_) );
NOR2_X1 U15525 ( .A1(n21113), .A2(n21110), .ZN(n21112) );
AND2_X1 U15526 ( .A1(n21113), .A2(n21110), .ZN(n21111) );
NAND2_X1 U15527 ( .A1(n21109), .A2(n21108), .ZN(n21110) );
NOR2_X1 U15528 ( .A1(n21153), .A2(n21152), .ZN(data_addr_o_20_) );
NOR2_X1 U15529 ( .A1(n21154), .A2(n21151), .ZN(n21153) );
AND2_X1 U15530 ( .A1(n21154), .A2(n21151), .ZN(n21152) );
NAND2_X1 U15531 ( .A1(n21150), .A2(n21149), .ZN(n21151) );
NOR2_X1 U15532 ( .A1(n21130), .A2(n21129), .ZN(data_addr_o_18_) );
NOR2_X1 U15533 ( .A1(n21136), .A2(n21128), .ZN(n21130) );
AND2_X1 U15534 ( .A1(n21136), .A2(n21128), .ZN(n21129) );
NAND2_X1 U15535 ( .A1(n21127), .A2(n21126), .ZN(n21128) );
NOR2_X1 U15536 ( .A1(n21103), .A2(n21102), .ZN(data_addr_o_15_) );
NOR2_X1 U15537 ( .A1(n21104), .A2(n21101), .ZN(n21103) );
AND2_X1 U15538 ( .A1(n21104), .A2(n21101), .ZN(n21102) );
NAND2_X1 U15539 ( .A1(n21100), .A2(n21099), .ZN(n21101) );
NOR2_X1 U15540 ( .A1(n21121), .A2(n21120), .ZN(data_addr_o_17_) );
AND2_X1 U15541 ( .A1(n21122), .A2(n21119), .ZN(n21120) );
NOR2_X1 U15542 ( .A1(n21122), .A2(n21119), .ZN(n21121) );
NAND2_X1 U15543 ( .A1(n21118), .A2(n21117), .ZN(n21119) );
NOR2_X1 U15544 ( .A1(n21144), .A2(n21143), .ZN(data_addr_o_19_) );
AND2_X1 U15545 ( .A1(n21145), .A2(n21142), .ZN(n21143) );
NOR2_X1 U15546 ( .A1(n21145), .A2(n21142), .ZN(n21144) );
NAND2_X1 U15547 ( .A1(n21141), .A2(n21140), .ZN(n21142) );
NOR2_X1 U15548 ( .A1(alu_adder_result_ex_1), .A2(data_addr_o_19_), .ZN(n21641) );
NOR2_X1 U15549 ( .A1(n21094), .A2(n21093), .ZN(data_addr_o_14_) );
NOR2_X1 U15550 ( .A1(n21095), .A2(n21092), .ZN(n21094) );
AND2_X1 U15551 ( .A1(n21095), .A2(n21092), .ZN(n21093) );
NAND2_X1 U15552 ( .A1(n21091), .A2(n21090), .ZN(n21092) );
NOR2_X1 U15553 ( .A1(n21085), .A2(n21084), .ZN(data_addr_o_13_) );
NOR2_X1 U15554 ( .A1(n21086), .A2(n21083), .ZN(n21085) );
AND2_X1 U15555 ( .A1(n21086), .A2(n21083), .ZN(n21084) );
NAND2_X1 U15556 ( .A1(n21082), .A2(n21081), .ZN(n21083) );
INV_X1 U15557 ( .A(data_addr_o_12_), .ZN(n20700) );
NOR2_X1 U15558 ( .A1(data_addr_o_9_), .A2(data_addr_o_8_), .ZN(n21625) );
NAND2_X1 U15559 ( .A1(n21636), .A2(n21635), .ZN(n21637) );
NOR2_X1 U15560 ( .A1(data_addr_o_10_), .A2(alu_adder_result_ex_0), .ZN(n21636) );
NOR2_X1 U15561 ( .A1(data_addr_o_12_), .A2(data_addr_o_11_), .ZN(n21635) );
INV_X1 U15562 ( .A(n92), .ZN(n20820) );
NAND2_X1 U15563 ( .A1(n1413), .A2(n20961), .ZN(n1318) );
NAND2_X1 U15564 ( .A1(n386), .A2(n359), .ZN(n1334) );
INV_X1 U15565 ( .A(n9927), .ZN(n20868) );
INV_X1 U15566 ( .A(data_addr_o_8_), .ZN(n20716) );
INV_X1 U15567 ( .A(data_addr_o_6_), .ZN(n20727) );
INV_X1 U15568 ( .A(data_addr_o_9_), .ZN(n20712) );
INV_X1 U15569 ( .A(data_addr_o_7_), .ZN(n20721) );
INV_X1 U15570 ( .A(data_addr_o_10_), .ZN(n20708) );
INV_X1 U15571 ( .A(n8104), .ZN(n16384) );
NAND2_X1 U15572 ( .A1(n7033), .A2(n9984), .ZN(n8624) );
INV_X1 U15573 ( .A(data_addr_o_11_), .ZN(n20704) );
NOR2_X1 U15574 ( .A1(data_addr_o_5_), .A2(data_addr_o_4_), .ZN(n21627) );
AND2_X1 U15575 ( .A1(n20868), .A2(n9984), .ZN(n16201) );
AND2_X1 U15576 ( .A1(n1413), .A2(n1423), .ZN(n1419) );
NAND2_X1 U15577 ( .A1(n9909), .A2(n20852), .ZN(n8575) );
NOR2_X1 U15578 ( .A1(n9908), .A2(n20823), .ZN(n9909) );
NAND2_X1 U15579 ( .A1(n9789), .A2(n20858), .ZN(n8685) );
BUF_X1 U15580 ( .A(n8584), .Z(n16372) );
BUF_X1 U15581 ( .A(n8567), .Z(n16375) );
AND2_X1 U15582 ( .A1(n21706), .A2(n20863), .ZN(n22081) );
BUF_X1 U15583 ( .A(n78), .Z(n16471) );
BUF_X1 U15584 ( .A(n22011), .Z(n16358) );
BUF_X1 U15585 ( .A(n8572), .Z(n16374) );
INV_X1 U15586 ( .A(n22009), .ZN(n20848) );
NOR2_X1 U15587 ( .A1(n21929), .A2(n20863), .ZN(n21951) );
INV_X1 U15588 ( .A(n8677), .ZN(n20826) );
NOR2_X1 U15589 ( .A1(n8121), .A2(n9918), .ZN(n9868) );
NOR2_X1 U15590 ( .A1(n20843), .A2(n8101), .ZN(n9907) );
NAND2_X1 U15591 ( .A1(n20852), .A2(n20825), .ZN(n8688) );
INV_X1 U15592 ( .A(alu_adder_result_ex_1), .ZN(n20753) );
NAND2_X1 U15593 ( .A1(n9926), .A2(n9868), .ZN(n8751) );
NOR2_X1 U15594 ( .A1(n8115), .A2(n9927), .ZN(n9926) );
INV_X1 U15595 ( .A(alu_adder_result_ex_0), .ZN(n20757) );
NOR2_X1 U15596 ( .A1(n20824), .A2(n15796), .ZN(n8621) );
INV_X1 U15597 ( .A(n9362), .ZN(n20824) );
NAND2_X1 U15598 ( .A1(n21999), .A2(n21873), .ZN(ex_block_i_alu_i_shift_result_ext_signed_16) );
NAND2_X1 U15599 ( .A1(n21872), .A2(n20850), .ZN(n21873) );
NAND2_X1 U15600 ( .A1(n21999), .A2(n21881), .ZN(ex_block_i_alu_i_shift_result_ext_signed_17) );
NAND2_X1 U15601 ( .A1(n21907), .A2(n20850), .ZN(n21881) );
NAND2_X1 U15602 ( .A1(n21999), .A2(n21890), .ZN(ex_block_i_alu_i_shift_result_ext_signed_18) );
NAND2_X1 U15603 ( .A1(n21980), .A2(n20850), .ZN(n21890) );
NAND2_X1 U15604 ( .A1(n21999), .A2(n21900), .ZN(ex_block_i_alu_i_shift_result_ext_signed_19) );
NAND2_X1 U15605 ( .A1(n22006), .A2(n20850), .ZN(n21900) );
NAND2_X1 U15606 ( .A1(n21999), .A2(n21933), .ZN(ex_block_i_alu_i_shift_result_ext_signed_20) );
NAND2_X1 U15607 ( .A1(n22026), .A2(n20850), .ZN(n21933) );
NAND2_X1 U15608 ( .A1(n21999), .A2(n21939), .ZN(ex_block_i_alu_i_shift_result_ext_signed_21) );
NAND2_X1 U15609 ( .A1(n22036), .A2(n20850), .ZN(n21939) );
NAND2_X1 U15610 ( .A1(n21999), .A2(n21945), .ZN(ex_block_i_alu_i_shift_result_ext_signed_22) );
NAND2_X1 U15611 ( .A1(n22046), .A2(n20850), .ZN(n21945) );
NAND2_X1 U15612 ( .A1(n21999), .A2(n21954), .ZN(ex_block_i_alu_i_shift_result_ext_signed_23) );
NAND2_X1 U15613 ( .A1(n22056), .A2(n20850), .ZN(n21954) );
NAND2_X1 U15614 ( .A1(n21999), .A2(n21959), .ZN(ex_block_i_alu_i_shift_result_ext_signed_24) );
NAND2_X1 U15615 ( .A1(n22065), .A2(n20850), .ZN(n21959) );
NAND2_X1 U15616 ( .A1(n21999), .A2(n21965), .ZN(ex_block_i_alu_i_shift_result_ext_signed_25) );
NAND2_X1 U15617 ( .A1(n22075), .A2(n20850), .ZN(n21965) );
NAND2_X1 U15618 ( .A1(n21999), .A2(n21967), .ZN(ex_block_i_alu_i_shift_result_ext_signed_26) );
NAND2_X1 U15619 ( .A1(n21966), .A2(n20850), .ZN(n21967) );
NAND2_X1 U15620 ( .A1(n21999), .A2(n21969), .ZN(ex_block_i_alu_i_shift_result_ext_signed_27) );
NAND2_X1 U15621 ( .A1(n21968), .A2(n20850), .ZN(n21969) );
NAND2_X1 U15622 ( .A1(n21999), .A2(n21971), .ZN(ex_block_i_alu_i_shift_result_ext_signed_28) );
NAND2_X1 U15623 ( .A1(n21970), .A2(n20850), .ZN(n21971) );
NAND2_X1 U15624 ( .A1(n21999), .A2(n21973), .ZN(ex_block_i_alu_i_shift_result_ext_signed_29) );
NAND2_X1 U15625 ( .A1(n21972), .A2(n20850), .ZN(n21973) );
NAND2_X1 U15626 ( .A1(n21999), .A2(n21996), .ZN(ex_block_i_alu_i_shift_result_ext_signed_30) );
NAND2_X1 U15627 ( .A1(n21995), .A2(n20850), .ZN(n21996) );
INV_X1 U15628 ( .A(n8102), .ZN(n16386) );
INV_X1 U15629 ( .A(n21929), .ZN(n20130) );
NOR2_X1 U15630 ( .A1(n22055), .A2(n22074), .ZN(n22058) );
NOR2_X1 U15631 ( .A1(n22045), .A2(n22074), .ZN(n22048) );
NOR2_X1 U15632 ( .A1(n22035), .A2(n22074), .ZN(n22038) );
NOR2_X1 U15633 ( .A1(n22025), .A2(n22074), .ZN(n22028) );
NOR2_X1 U15634 ( .A1(n16359), .A2(n20134), .ZN(n21827) );
INV_X1 U15635 ( .A(data_addr_o_4_), .ZN(n20738) );
INV_X1 U15636 ( .A(data_addr_o_2_), .ZN(n20749) );
INV_X1 U15637 ( .A(data_addr_o_5_), .ZN(n20732) );
INV_X1 U15638 ( .A(data_addr_o_3_), .ZN(n20743) );
NOR2_X1 U15639 ( .A1(n20173), .A2(n21960), .ZN(n21948) );
NOR2_X1 U15640 ( .A1(n22025), .A2(n22078), .ZN(n21699) );
NOR2_X1 U15641 ( .A1(n20485), .A2(n22078), .ZN(n21871) );
NOR2_X1 U15642 ( .A1(n20524), .A2(n22078), .ZN(n21862) );
NOR2_X1 U15643 ( .A1(n20564), .A2(n22078), .ZN(n21854) );
NOR2_X1 U15644 ( .A1(n20604), .A2(n22078), .ZN(n21817) );
NOR2_X1 U15645 ( .A1(n20642), .A2(n22078), .ZN(n21808) );
NOR2_X1 U15646 ( .A1(n20677), .A2(n22078), .ZN(n21766) );
NOR2_X1 U15647 ( .A1(n20643), .A2(n22078), .ZN(n22085) );
NOR2_X1 U15648 ( .A1(n20605), .A2(n22078), .ZN(n22073) );
NOR2_X1 U15649 ( .A1(n20565), .A2(n22078), .ZN(n22064) );
NOR2_X1 U15650 ( .A1(n20525), .A2(n22078), .ZN(n22054) );
NOR2_X1 U15651 ( .A1(n20484), .A2(n22078), .ZN(n22044) );
NOR2_X1 U15652 ( .A1(n20444), .A2(n22078), .ZN(n22034) );
NOR2_X1 U15653 ( .A1(n22055), .A2(n22078), .ZN(n22008) );
NOR2_X1 U15654 ( .A1(n22045), .A2(n22078), .ZN(n21982) );
NOR2_X1 U15655 ( .A1(n22035), .A2(n22078), .ZN(n21909) );
INV_X1 U15656 ( .A(n9844), .ZN(n20852) );
NOR2_X1 U15657 ( .A1(n20288), .A2(n21949), .ZN(n21694) );
NOR2_X1 U15658 ( .A1(n20129), .A2(n21949), .ZN(n21942) );
NOR2_X1 U15659 ( .A1(n20131), .A2(n21949), .ZN(n21936) );
NOR2_X1 U15660 ( .A1(n20133), .A2(n21949), .ZN(n21930) );
NOR2_X1 U15661 ( .A1(n20173), .A2(n21949), .ZN(n21896) );
NOR2_X1 U15662 ( .A1(n20211), .A2(n21949), .ZN(n21886) );
NOR2_X1 U15663 ( .A1(n20249), .A2(n21949), .ZN(n21877) );
NAND2_X1 U15664 ( .A1(n21997), .A2(n20850), .ZN(n21998) );
NOR2_X1 U15665 ( .A1(n9925), .A2(n8118), .ZN(n9923) );
NAND2_X1 U15666 ( .A1(n16361), .A2(n9362), .ZN(n8945) );
NAND2_X1 U15667 ( .A1(n21860), .A2(n21859), .ZN(n21861) );
NAND2_X1 U15668 ( .A1(n20848), .A2(n21885), .ZN(n21860) );
NAND2_X1 U15669 ( .A1(n22081), .A2(n21882), .ZN(n21859) );
NAND2_X1 U15670 ( .A1(n21852), .A2(n21851), .ZN(n21853) );
NAND2_X1 U15671 ( .A1(n20848), .A2(n21962), .ZN(n21852) );
NAND2_X1 U15672 ( .A1(n22081), .A2(n22079), .ZN(n21851) );
NAND2_X1 U15673 ( .A1(n22083), .A2(n22082), .ZN(n22084) );
NAND2_X1 U15674 ( .A1(n20848), .A2(n22079), .ZN(n22083) );
NAND2_X1 U15675 ( .A1(n22081), .A2(n22080), .ZN(n22082) );
NOR2_X1 U15676 ( .A1(n20605), .A2(n22009), .ZN(n21723) );
NOR2_X1 U15677 ( .A1(n20642), .A2(n22009), .ZN(n22024) );
NOR2_X1 U15678 ( .A1(n20677), .A2(n22009), .ZN(n21994) );
NOR2_X1 U15679 ( .A1(n20643), .A2(n22009), .ZN(n21926) );
NOR2_X1 U15680 ( .A1(n20135), .A2(n15801), .ZN(n384) );
NOR2_X1 U15681 ( .A1(n20128), .A2(n21894), .ZN(n21897) );
NOR2_X1 U15682 ( .A1(n20129), .A2(n21894), .ZN(n21887) );
NOR2_X1 U15683 ( .A1(n20133), .A2(n21894), .ZN(n21695) );
NOR2_X1 U15684 ( .A1(n20131), .A2(n21894), .ZN(n21878) );
NOR2_X1 U15685 ( .A1(n20845), .A2(n20827), .ZN(n9989) );
NAND2_X1 U15686 ( .A1(n21944), .A2(n21943), .ZN(n22046) );
NOR2_X1 U15687 ( .A1(n21941), .A2(n21940), .ZN(n21944) );
NOR2_X1 U15688 ( .A1(n21951), .A2(n21942), .ZN(n21943) );
NOR2_X1 U15689 ( .A1(n20211), .A2(n21960), .ZN(n21941) );
NAND2_X1 U15690 ( .A1(n21938), .A2(n21937), .ZN(n22036) );
NOR2_X1 U15691 ( .A1(n21935), .A2(n21934), .ZN(n21938) );
NOR2_X1 U15692 ( .A1(n21951), .A2(n21936), .ZN(n21937) );
NOR2_X1 U15693 ( .A1(n20249), .A2(n21960), .ZN(n21935) );
INV_X1 U15694 ( .A(n21855), .ZN(n20129) );
INV_X1 U15695 ( .A(n22030), .ZN(n20605) );
INV_X1 U15696 ( .A(n22060), .ZN(n20642) );
INV_X1 U15697 ( .A(n22050), .ZN(n20677) );
INV_X1 U15698 ( .A(n22040), .ZN(n20643) );
INV_X1 U15699 ( .A(n21863), .ZN(n20128) );
NAND2_X1 U15700 ( .A1(alu_adder_result_ex_0), .A2(n20753), .ZN(n6318) );
INV_X1 U15701 ( .A(n9918), .ZN(n20860) );
NAND2_X1 U15702 ( .A1(n9938), .A2(n20868), .ZN(n8591) );
NAND2_X1 U15703 ( .A1(n9938), .A2(n7033), .ZN(n8585) );
NAND2_X1 U15704 ( .A1(n20827), .A2(n9973), .ZN(n10034) );
NAND2_X1 U15705 ( .A1(n21687), .A2(n21686), .ZN(n21810) );
NOR2_X1 U15706 ( .A1(n21685), .A2(n21684), .ZN(n21686) );
NOR2_X1 U15707 ( .A1(n21683), .A2(n21682), .ZN(n21687) );
NOR2_X1 U15708 ( .A1(n22015), .A2(n20134), .ZN(n21684) );
NAND2_X1 U15709 ( .A1(n21829), .A2(n21828), .ZN(n21876) );
NOR2_X1 U15710 ( .A1(n21827), .A2(n21826), .ZN(n21828) );
NOR2_X1 U15711 ( .A1(n21825), .A2(n21824), .ZN(n21829) );
NOR2_X1 U15712 ( .A1(n22015), .A2(n20132), .ZN(n21826) );
INV_X1 U15713 ( .A(n8122), .ZN(n20832) );
INV_X1 U15714 ( .A(ex_block_i_alu_i_N294), .ZN(n20132) );
NAND2_X1 U15715 ( .A1(n21865), .A2(n21864), .ZN(n21997) );
NAND2_X1 U15716 ( .A1(n20855), .A2(n21863), .ZN(n21864) );
INV_X1 U15717 ( .A(n9908), .ZN(n20837) );
NAND2_X1 U15718 ( .A1(n21865), .A2(n21856), .ZN(n21995) );
NAND2_X1 U15719 ( .A1(n20855), .A2(n21855), .ZN(n21856) );
NAND2_X1 U15720 ( .A1(n21865), .A2(n21830), .ZN(n21972) );
NAND2_X1 U15721 ( .A1(n20855), .A2(n21876), .ZN(n21830) );
NAND2_X1 U15722 ( .A1(n21865), .A2(n21811), .ZN(n21970) );
NAND2_X1 U15723 ( .A1(n20855), .A2(n21810), .ZN(n21811) );
NAND2_X1 U15724 ( .A1(n21784), .A2(n21783), .ZN(n21968) );
NAND2_X1 U15725 ( .A1(n20855), .A2(n21895), .ZN(n21783) );
NOR2_X1 U15726 ( .A1(n20130), .A2(n21776), .ZN(n21784) );
NOR2_X1 U15727 ( .A1(n20128), .A2(n21960), .ZN(n21776) );
NAND2_X1 U15728 ( .A1(n21742), .A2(n21741), .ZN(n21966) );
NAND2_X1 U15729 ( .A1(n20855), .A2(n21885), .ZN(n21741) );
NOR2_X1 U15730 ( .A1(n20130), .A2(n21734), .ZN(n21742) );
NOR2_X1 U15731 ( .A1(n20129), .A2(n21960), .ZN(n21734) );
NAND2_X1 U15732 ( .A1(n21964), .A2(n21963), .ZN(n22075) );
NAND2_X1 U15733 ( .A1(n20855), .A2(n21962), .ZN(n21963) );
NOR2_X1 U15734 ( .A1(n20130), .A2(n21961), .ZN(n21964) );
NOR2_X1 U15735 ( .A1(n20131), .A2(n21960), .ZN(n21961) );
NAND2_X1 U15736 ( .A1(n21958), .A2(n21957), .ZN(n22065) );
NAND2_X1 U15737 ( .A1(n20855), .A2(n21956), .ZN(n21957) );
NOR2_X1 U15738 ( .A1(n20130), .A2(n21955), .ZN(n21958) );
NOR2_X1 U15739 ( .A1(n20133), .A2(n21960), .ZN(n21955) );
INV_X1 U15740 ( .A(n22069), .ZN(n20604) );
INV_X1 U15741 ( .A(n22068), .ZN(n20445) );
INV_X1 U15742 ( .A(n21956), .ZN(n20288) );
INV_X1 U15743 ( .A(n22059), .ZN(n20485) );
INV_X1 U15744 ( .A(n22049), .ZN(n20524) );
INV_X1 U15745 ( .A(n21895), .ZN(n20173) );
INV_X1 U15746 ( .A(n21891), .ZN(n20327) );
INV_X1 U15747 ( .A(n21885), .ZN(n20211) );
INV_X1 U15748 ( .A(n21882), .ZN(n20366) );
INV_X1 U15749 ( .A(n21962), .ZN(n20249) );
INV_X1 U15750 ( .A(n22080), .ZN(n20564) );
INV_X1 U15751 ( .A(n22079), .ZN(n20405) );
NAND2_X1 U15752 ( .A1(n21953), .A2(n21952), .ZN(n22056) );
NOR2_X1 U15753 ( .A1(n21951), .A2(n21950), .ZN(n21952) );
NOR2_X1 U15754 ( .A1(n21948), .A2(n21947), .ZN(n21953) );
NOR2_X1 U15755 ( .A1(n20128), .A2(n21949), .ZN(n21950) );
NAND2_X1 U15756 ( .A1(n21932), .A2(n21931), .ZN(n22026) );
NOR2_X1 U15757 ( .A1(n21928), .A2(n21927), .ZN(n21932) );
NOR2_X1 U15758 ( .A1(n21951), .A2(n21930), .ZN(n21931) );
NOR2_X1 U15759 ( .A1(n20288), .A2(n21960), .ZN(n21928) );
INV_X1 U15760 ( .A(n9925), .ZN(n20844) );
INV_X1 U15761 ( .A(n22029), .ZN(n20444) );
INV_X1 U15762 ( .A(n22010), .ZN(n20565) );
INV_X1 U15763 ( .A(n21983), .ZN(n20525) );
INV_X1 U15764 ( .A(n22039), .ZN(n20484) );
NAND2_X1 U15765 ( .A1(n9913), .A2(n20852), .ZN(n8576) );
NOR2_X1 U15766 ( .A1(n9841), .A2(n20823), .ZN(n9913) );
NAND2_X1 U15767 ( .A1(n21697), .A2(n21696), .ZN(n21872) );
NOR2_X1 U15768 ( .A1(n21681), .A2(n21680), .ZN(n21697) );
NOR2_X1 U15769 ( .A1(n21695), .A2(n21694), .ZN(n21696) );
NOR2_X1 U15770 ( .A1(n20445), .A2(n21960), .ZN(n21681) );
NAND2_X1 U15771 ( .A1(n21899), .A2(n21898), .ZN(n22006) );
NOR2_X1 U15772 ( .A1(n21893), .A2(n21892), .ZN(n21899) );
NOR2_X1 U15773 ( .A1(n21897), .A2(n21896), .ZN(n21898) );
NOR2_X1 U15774 ( .A1(n20327), .A2(n21960), .ZN(n21893) );
NAND2_X1 U15775 ( .A1(n21889), .A2(n21888), .ZN(n21980) );
NOR2_X1 U15776 ( .A1(n21884), .A2(n21883), .ZN(n21889) );
NOR2_X1 U15777 ( .A1(n21887), .A2(n21886), .ZN(n21888) );
NOR2_X1 U15778 ( .A1(n20366), .A2(n21960), .ZN(n21884) );
NAND2_X1 U15779 ( .A1(n21880), .A2(n21879), .ZN(n21907) );
NOR2_X1 U15780 ( .A1(n21875), .A2(n21874), .ZN(n21880) );
NOR2_X1 U15781 ( .A1(n21878), .A2(n21877), .ZN(n21879) );
NOR2_X1 U15782 ( .A1(n20405), .A2(n21960), .ZN(n21875) );
INV_X1 U15783 ( .A(n7311), .ZN(n20858) );
NAND2_X1 U15784 ( .A1(n9789), .A2(n20857), .ZN(n8590) );
INV_X1 U15785 ( .A(n6697), .ZN(n20857) );
NOR2_X1 U15786 ( .A1(n16203), .A2(n16204), .ZN(n16202) );
OR2_X1 U15787 ( .A1(n22008), .A2(n22007), .ZN(n16203) );
OR2_X1 U15788 ( .A1(n22024), .A2(n22023), .ZN(n16204) );
NOR2_X1 U15789 ( .A1(n16206), .A2(n16207), .ZN(n16205) );
OR2_X1 U15790 ( .A1(n21982), .A2(n21981), .ZN(n16206) );
OR2_X1 U15791 ( .A1(n21994), .A2(n21993), .ZN(n16207) );
NOR2_X1 U15792 ( .A1(n16209), .A2(n16210), .ZN(n16208) );
OR2_X1 U15793 ( .A1(n21909), .A2(n21908), .ZN(n16209) );
OR2_X1 U15794 ( .A1(n21926), .A2(n21925), .ZN(n16210) );
NOR2_X1 U15795 ( .A1(n16212), .A2(n16213), .ZN(n16211) );
OR2_X1 U15796 ( .A1(n21813), .A2(n21812), .ZN(n16212) );
OR2_X1 U15797 ( .A1(n21817), .A2(n21816), .ZN(n16213) );
NOR2_X1 U15798 ( .A1(n16215), .A2(n16216), .ZN(n16214) );
OR2_X1 U15799 ( .A1(n21786), .A2(n21785), .ZN(n16215) );
OR2_X1 U15800 ( .A1(n21808), .A2(n21807), .ZN(n16216) );
NOR2_X1 U15801 ( .A1(n16218), .A2(n16219), .ZN(n16217) );
OR2_X1 U15802 ( .A1(n22067), .A2(n22066), .ZN(n16218) );
OR2_X1 U15803 ( .A1(n22073), .A2(n22072), .ZN(n16219) );
NOR2_X1 U15804 ( .A1(n16221), .A2(n16222), .ZN(n16220) );
OR2_X1 U15805 ( .A1(n22058), .A2(n22057), .ZN(n16221) );
OR2_X1 U15806 ( .A1(n22064), .A2(n22063), .ZN(n16222) );
NAND2_X1 U15807 ( .A1(n20837), .A2(n20827), .ZN(n9953) );
NAND2_X1 U15808 ( .A1(n21869), .A2(n21868), .ZN(n21870) );
NAND2_X1 U15809 ( .A1(n20848), .A2(n21895), .ZN(n21869) );
NAND2_X1 U15810 ( .A1(n22081), .A2(n21891), .ZN(n21868) );
NAND2_X1 U15811 ( .A1(n21815), .A2(n21814), .ZN(n21816) );
NAND2_X1 U15812 ( .A1(n20848), .A2(n21956), .ZN(n21815) );
NAND2_X1 U15813 ( .A1(n22081), .A2(n22068), .ZN(n21814) );
NAND2_X1 U15814 ( .A1(n21806), .A2(n21805), .ZN(n21807) );
NAND2_X1 U15815 ( .A1(n20848), .A2(n21891), .ZN(n21806) );
NAND2_X1 U15816 ( .A1(n22081), .A2(n22059), .ZN(n21805) );
NAND2_X1 U15817 ( .A1(n21764), .A2(n21763), .ZN(n21765) );
NAND2_X1 U15818 ( .A1(n20848), .A2(n21882), .ZN(n21764) );
NAND2_X1 U15819 ( .A1(n22081), .A2(n22049), .ZN(n21763) );
NAND2_X1 U15820 ( .A1(n22071), .A2(n22070), .ZN(n22072) );
NAND2_X1 U15821 ( .A1(n20848), .A2(n22068), .ZN(n22071) );
NAND2_X1 U15822 ( .A1(n22081), .A2(n22069), .ZN(n22070) );
NAND2_X1 U15823 ( .A1(n22062), .A2(n22061), .ZN(n22063) );
NAND2_X1 U15824 ( .A1(n22081), .A2(n22060), .ZN(n22061) );
NAND2_X1 U15825 ( .A1(n20848), .A2(n22059), .ZN(n22062) );
NAND2_X1 U15826 ( .A1(n22052), .A2(n22051), .ZN(n22053) );
NAND2_X1 U15827 ( .A1(n22081), .A2(n22050), .ZN(n22051) );
NAND2_X1 U15828 ( .A1(n20848), .A2(n22049), .ZN(n22052) );
NAND2_X1 U15829 ( .A1(n22042), .A2(n22041), .ZN(n22043) );
NAND2_X1 U15830 ( .A1(n22081), .A2(n22040), .ZN(n22041) );
NAND2_X1 U15831 ( .A1(n20848), .A2(n22080), .ZN(n22042) );
NAND2_X1 U15832 ( .A1(n22032), .A2(n22031), .ZN(n22033) );
NAND2_X1 U15833 ( .A1(n22081), .A2(n22030), .ZN(n22031) );
NAND2_X1 U15834 ( .A1(n20848), .A2(n22069), .ZN(n22032) );
NAND2_X1 U15835 ( .A1(n21721), .A2(n21720), .ZN(n21722) );
NAND2_X1 U15836 ( .A1(n22081), .A2(n22029), .ZN(n21721) );
NAND2_X1 U15837 ( .A1(n20849), .A2(n21719), .ZN(n21720) );
NAND2_X1 U15838 ( .A1(n21718), .A2(n21717), .ZN(n21719) );
NAND2_X1 U15839 ( .A1(n22022), .A2(n22021), .ZN(n22023) );
NAND2_X1 U15840 ( .A1(n22081), .A2(n22010), .ZN(n22022) );
NAND2_X1 U15841 ( .A1(n20849), .A2(n22020), .ZN(n22021) );
NAND2_X1 U15842 ( .A1(n22019), .A2(n22018), .ZN(n22020) );
NAND2_X1 U15843 ( .A1(n21992), .A2(n21991), .ZN(n21993) );
NAND2_X1 U15844 ( .A1(n22081), .A2(n21983), .ZN(n21992) );
NAND2_X1 U15845 ( .A1(n20849), .A2(n21990), .ZN(n21991) );
NAND2_X1 U15846 ( .A1(n21989), .A2(n21988), .ZN(n21990) );
NAND2_X1 U15847 ( .A1(n21924), .A2(n21923), .ZN(n21925) );
NAND2_X1 U15848 ( .A1(n22081), .A2(n22039), .ZN(n21924) );
NAND2_X1 U15849 ( .A1(n20849), .A2(n21922), .ZN(n21923) );
NAND2_X1 U15850 ( .A1(n21921), .A2(n21920), .ZN(n21922) );
NOR2_X1 U15851 ( .A1(n16224), .A2(n16225), .ZN(n16223) );
OR2_X1 U15852 ( .A1(n21867), .A2(n21866), .ZN(n16224) );
OR2_X1 U15853 ( .A1(n21871), .A2(n21870), .ZN(n16225) );
NOR2_X1 U15854 ( .A1(n16227), .A2(n16228), .ZN(n16226) );
OR2_X1 U15855 ( .A1(n21858), .A2(n21857), .ZN(n16227) );
OR2_X1 U15856 ( .A1(n21862), .A2(n21861), .ZN(n16228) );
NOR2_X1 U15857 ( .A1(n16230), .A2(n16231), .ZN(n16229) );
OR2_X1 U15858 ( .A1(n21832), .A2(n21831), .ZN(n16230) );
OR2_X1 U15859 ( .A1(n21854), .A2(n21853), .ZN(n16231) );
NOR2_X1 U15860 ( .A1(n16233), .A2(n16234), .ZN(n16232) );
OR2_X1 U15861 ( .A1(n21744), .A2(n21743), .ZN(n16233) );
OR2_X1 U15862 ( .A1(n21766), .A2(n21765), .ZN(n16234) );
NOR2_X1 U15863 ( .A1(n16236), .A2(n16237), .ZN(n16235) );
OR2_X1 U15864 ( .A1(n22077), .A2(n22076), .ZN(n16236) );
OR2_X1 U15865 ( .A1(n22085), .A2(n22084), .ZN(n16237) );
NOR2_X1 U15866 ( .A1(n16239), .A2(n16240), .ZN(n16238) );
OR2_X1 U15867 ( .A1(n22048), .A2(n22047), .ZN(n16239) );
OR2_X1 U15868 ( .A1(n22054), .A2(n22053), .ZN(n16240) );
NOR2_X1 U15869 ( .A1(n16242), .A2(n16243), .ZN(n16241) );
OR2_X1 U15870 ( .A1(n22038), .A2(n22037), .ZN(n16242) );
OR2_X1 U15871 ( .A1(n22044), .A2(n22043), .ZN(n16243) );
NOR2_X1 U15872 ( .A1(n16245), .A2(n16246), .ZN(n16244) );
OR2_X1 U15873 ( .A1(n22028), .A2(n22027), .ZN(n16245) );
OR2_X1 U15874 ( .A1(n22034), .A2(n22033), .ZN(n16246) );
NOR2_X1 U15875 ( .A1(n16248), .A2(n16249), .ZN(n16247) );
OR2_X1 U15876 ( .A1(n21699), .A2(n21698), .ZN(n16248) );
OR2_X1 U15877 ( .A1(n21723), .A2(n21722), .ZN(n16249) );
INV_X1 U15878 ( .A(n21773), .ZN(n20866) );
BUF_X1 U15879 ( .A(n19966), .Z(n16346) );
INV_X1 U15880 ( .A(n8083), .ZN(n19969) );
INV_X1 U15881 ( .A(n8773), .ZN(n20947) );
NAND2_X1 U15882 ( .A1(n7310), .A2(n19983), .ZN(n7257) );
NOR2_X1 U15883 ( .A1(n7311), .A2(n6698), .ZN(n7310) );
INV_X1 U15884 ( .A(n3776), .ZN(n20925) );
BUF_X1 U15885 ( .A(n7323), .Z(n16392) );
BUF_X1 U15886 ( .A(n4066), .Z(n16426) );
BUF_X1 U15887 ( .A(n5385), .Z(n16414) );
BUF_X1 U15888 ( .A(n8456), .Z(n16377) );
INV_X1 U15889 ( .A(n6711), .ZN(n19974) );
INV_X1 U15890 ( .A(n4797), .ZN(n20907) );
BUF_X1 U15891 ( .A(n5382), .Z(n16415) );
BUF_X1 U15892 ( .A(n5278), .Z(n16416) );
BUF_X1 U15893 ( .A(n5277), .Z(n16417) );
INV_X1 U15894 ( .A(n5904), .ZN(n20939) );
BUF_X1 U15895 ( .A(n7876), .Z(n16387) );
NOR2_X1 U15896 ( .A1(n4046), .A2(n4005), .ZN(n3773) );
NOR2_X1 U15897 ( .A1(n20928), .A2(n4005), .ZN(n3774) );
BUF_X1 U15898 ( .A(n20950), .Z(n16356) );
BUF_X1 U15899 ( .A(n4280), .Z(n16422) );
NAND2_X1 U15900 ( .A1(n16404), .A2(n6694), .ZN(n6561) );
NAND2_X1 U15901 ( .A1(n6695), .A2(n19983), .ZN(n6694) );
NOR2_X1 U15902 ( .A1(n6697), .A2(n6698), .ZN(n6695) );
BUF_X1 U15903 ( .A(n5826), .Z(n16409) );
BUF_X1 U15904 ( .A(n20961), .Z(n16357) );
BUF_X1 U15905 ( .A(n7319), .Z(n16395) );
BUF_X1 U15906 ( .A(n20023), .Z(n16350) );
INV_X1 U15907 ( .A(n5911), .ZN(n20958) );
BUF_X1 U15908 ( .A(n8601), .Z(n16364) );
BUF_X1 U15909 ( .A(n20931), .Z(n16355) );
BUF_X1 U15910 ( .A(n6719), .Z(n16402) );
INV_X1 U15911 ( .A(n16461), .ZN(n16460) );
BUF_X1 U15912 ( .A(n5818), .Z(n16410) );
INV_X1 U15913 ( .A(n1452), .ZN(n16465) );
INV_X1 U15914 ( .A(n15811), .ZN(n16412) );
INV_X1 U15915 ( .A(n15811), .ZN(n16411) );
NAND2_X1 U15916 ( .A1(n16450), .A2(n2704), .ZN(n2117) );
NAND2_X1 U15917 ( .A1(n19901), .A2(n19903), .ZN(n2704) );
INV_X1 U15918 ( .A(n2142), .ZN(n19881) );
AND2_X1 U15919 ( .A1(n5910), .A2(n6186), .ZN(n6079) );
INV_X1 U15920 ( .A(n7226), .ZN(n19809) );
NOR2_X1 U15921 ( .A1(n19940), .A2(n19894), .ZN(n2025) );
NAND2_X1 U15922 ( .A1(n19909), .A2(n2142), .ZN(n2036) );
INV_X1 U15923 ( .A(n7037), .ZN(n19805) );
OR2_X1 U15924 ( .A1(n7716), .A2(n7717), .ZN(n7562) );
NAND2_X1 U15925 ( .A1(n7795), .A2(n19983), .ZN(n7725) );
INV_X1 U15926 ( .A(n7194), .ZN(n19803) );
BUF_X1 U15927 ( .A(n8436), .Z(n16379) );
NAND2_X1 U15928 ( .A1(n10157), .A2(n10158), .ZN(n10022) );
BUF_X1 U15929 ( .A(n3740), .Z(n16428) );
NAND2_X1 U15930 ( .A1(n7076), .A2(n7077), .ZN(n7040) );
NAND2_X1 U15931 ( .A1(n7078), .A2(n19983), .ZN(n7077) );
NOR2_X1 U15932 ( .A1(n16400), .A2(n20929), .ZN(n7076) );
INV_X1 U15933 ( .A(n7577), .ZN(n19975) );
NAND2_X1 U15934 ( .A1(n19983), .A2(n16386), .ZN(n7803) );
NAND2_X1 U15935 ( .A1(n2332), .A2(n2142), .ZN(n2109) );
INV_X1 U15936 ( .A(n7041), .ZN(n20929) );
NOR2_X1 U15937 ( .A1(n10501), .A2(n20956), .ZN(n10505) );
BUF_X1 U15938 ( .A(n5904), .Z(n16334) );
INV_X1 U15939 ( .A(n2184), .ZN(n19894) );
NAND2_X1 U15940 ( .A1(n2675), .A2(n19906), .ZN(n2470) );
NAND2_X1 U15941 ( .A1(n19941), .A2(n19940), .ZN(n2696) );
NOR2_X1 U15942 ( .A1(n2180), .A2(n2233), .ZN(n2202) );
AND2_X1 U15943 ( .A1(n1885), .A2(n2234), .ZN(n2233) );
NAND2_X1 U15944 ( .A1(n2182), .A2(n2235), .ZN(n2234) );
NOR2_X1 U15945 ( .A1(n2025), .A2(n2026), .ZN(n2015) );
INV_X1 U15946 ( .A(n8306), .ZN(n19980) );
NOR2_X1 U15947 ( .A1(n20876), .A2(n4036), .ZN(n7612) );
INV_X1 U15948 ( .A(n2471), .ZN(n19876) );
NAND2_X1 U15949 ( .A1(n19983), .A2(n7040), .ZN(n7052) );
NAND2_X1 U15950 ( .A1(n9843), .A2(n19983), .ZN(n8883) );
NOR2_X1 U15951 ( .A1(n8101), .A2(n9844), .ZN(n9843) );
INV_X1 U15952 ( .A(n8079), .ZN(n19978) );
NOR2_X1 U15953 ( .A1(n2113), .A2(n19939), .ZN(n2649) );
AND2_X1 U15954 ( .A1(n9840), .A2(n19983), .ZN(n8310) );
NOR2_X1 U15955 ( .A1(n9841), .A2(n8121), .ZN(n9840) );
INV_X1 U15956 ( .A(n3567), .ZN(n19884) );
NOR2_X1 U15957 ( .A1(n19863), .A2(n2901), .ZN(n3013) );
NOR2_X1 U15958 ( .A1(n19851), .A2(n16443), .ZN(n2993) );
NOR2_X1 U15959 ( .A1(n19841), .A2(n2901), .ZN(n2977) );
NOR2_X1 U15960 ( .A1(n19828), .A2(n16443), .ZN(n2957) );
NOR2_X1 U15961 ( .A1(n19823), .A2(n2901), .ZN(n2949) );
NOR2_X1 U15962 ( .A1(n19821), .A2(n2901), .ZN(n2945) );
NAND2_X1 U15963 ( .A1(n20906), .A2(n20999), .ZN(n4061) );
NAND2_X1 U15964 ( .A1(n16451), .A2(n2059), .ZN(n2138) );
NOR2_X1 U15965 ( .A1(n8414), .A2(n19980), .ZN(n8149) );
NOR2_X1 U15966 ( .A1(alu_adder_result_ex_0), .A2(n4287), .ZN(n4727) );
NAND2_X1 U15967 ( .A1(n8119), .A2(n20825), .ZN(n6698) );
NOR2_X1 U15968 ( .A1(n8121), .A2(n8122), .ZN(n8119) );
NOR2_X1 U15969 ( .A1(n19749), .A2(n16378), .ZN(n8890) );
NOR2_X1 U15970 ( .A1(n19751), .A2(n16377), .ZN(n8459) );
NOR2_X1 U15971 ( .A1(n19755), .A2(n8169), .ZN(n8180) );
NOR2_X1 U15972 ( .A1(n20712), .A2(n5386), .ZN(n5383) );
NOR2_X1 U15973 ( .A1(n20716), .A2(n5386), .ZN(n5390) );
NOR2_X1 U15974 ( .A1(n20721), .A2(n5386), .ZN(n5395) );
NOR2_X1 U15975 ( .A1(n20727), .A2(n5386), .ZN(n5400) );
NOR2_X1 U15976 ( .A1(n20732), .A2(n5386), .ZN(n5404) );
NOR2_X1 U15977 ( .A1(n20738), .A2(n5386), .ZN(n5408) );
NOR2_X1 U15978 ( .A1(n20743), .A2(n5386), .ZN(n5413) );
NOR2_X1 U15979 ( .A1(n20112), .A2(n5386), .ZN(n5417) );
NOR2_X1 U15980 ( .A1(n19801), .A2(n16381), .ZN(n8184) );
NOR2_X1 U15981 ( .A1(n19749), .A2(n16381), .ZN(n8316) );
NOR2_X1 U15982 ( .A1(n19801), .A2(n16378), .ZN(n8471) );
NOR2_X1 U15983 ( .A1(n19757), .A2(n8169), .ZN(n8188) );
NOR2_X1 U15984 ( .A1(n19757), .A2(n16377), .ZN(n8475) );
NOR2_X1 U15985 ( .A1(n19759), .A2(n8169), .ZN(n8192) );
NOR2_X1 U15986 ( .A1(n19759), .A2(n16377), .ZN(n8479) );
NOR2_X1 U15987 ( .A1(n19761), .A2(n8169), .ZN(n8196) );
NOR2_X1 U15988 ( .A1(n19761), .A2(n16377), .ZN(n8483) );
NOR2_X1 U15989 ( .A1(n19763), .A2(n8169), .ZN(n8200) );
NOR2_X1 U15990 ( .A1(n19763), .A2(n16377), .ZN(n8487) );
NOR2_X1 U15991 ( .A1(n19793), .A2(n16381), .ZN(n8147) );
NOR2_X1 U15992 ( .A1(n19793), .A2(n16378), .ZN(n8434) );
NOR2_X1 U15993 ( .A1(n19795), .A2(n16381), .ZN(n8153) );
NOR2_X1 U15994 ( .A1(n19795), .A2(n16378), .ZN(n8440) );
NOR2_X1 U15995 ( .A1(n19799), .A2(n16381), .ZN(n8161) );
NOR2_X1 U15996 ( .A1(n19799), .A2(n16378), .ZN(n8448) );
NOR2_X1 U15997 ( .A1(n19797), .A2(n16381), .ZN(n8157) );
NOR2_X1 U15998 ( .A1(n19797), .A2(n16378), .ZN(n8444) );
NOR2_X1 U15999 ( .A1(n19755), .A2(n16377), .ZN(n8467) );
NOR2_X1 U16000 ( .A1(n19753), .A2(n8169), .ZN(n8176) );
NOR2_X1 U16001 ( .A1(n19751), .A2(n8169), .ZN(n8172) );
NOR2_X1 U16002 ( .A1(n19749), .A2(n8169), .ZN(n8166) );
NOR2_X1 U16003 ( .A1(n19753), .A2(n16377), .ZN(n8463) );
NOR2_X1 U16004 ( .A1(n19749), .A2(n16377), .ZN(n8453) );
NOR2_X1 U16005 ( .A1(n20753), .A2(n5386), .ZN(n5473) );
NAND2_X1 U16006 ( .A1(n6702), .A2(n6703), .ZN(n4046) );
NOR2_X1 U16007 ( .A1(n20929), .A2(n20991), .ZN(n6702) );
NOR2_X1 U16008 ( .A1(n20989), .A2(n20985), .ZN(n6703) );
NAND2_X1 U16009 ( .A1(n20931), .A2(n7041), .ZN(n7717) );
NAND2_X1 U16010 ( .A1(n2049), .A2(n16452), .ZN(n2457) );
NAND2_X1 U16011 ( .A1(n19894), .A2(n2356), .ZN(n2238) );
NOR2_X1 U16012 ( .A1(n16439), .A2(n19863), .ZN(n3547) );
NOR2_X1 U16013 ( .A1(n19789), .A2(n16391), .ZN(n8048) );
NOR2_X1 U16014 ( .A1(n19779), .A2(n16390), .ZN(n8018) );
NOR2_X1 U16015 ( .A1(n19781), .A2(n16391), .ZN(n8024) );
NOR2_X1 U16016 ( .A1(n19783), .A2(n16390), .ZN(n8030) );
NOR2_X1 U16017 ( .A1(n19785), .A2(n16391), .ZN(n8036) );
NOR2_X1 U16018 ( .A1(n19787), .A2(n16390), .ZN(n8042) );
NOR2_X1 U16019 ( .A1(n19791), .A2(n16391), .ZN(n8054) );
NOR2_X1 U16020 ( .A1(n19753), .A2(n8150), .ZN(n8328) );
NOR2_X1 U16021 ( .A1(n19811), .A2(n8150), .ZN(n8412) );
NOR2_X1 U16022 ( .A1(n19751), .A2(n8150), .ZN(n8320) );
NOR2_X1 U16023 ( .A1(n19807), .A2(n8150), .ZN(n8324) );
NOR2_X1 U16024 ( .A1(n19769), .A2(n8150), .ZN(n8360) );
NOR2_X1 U16025 ( .A1(n19751), .A2(n8437), .ZN(n8925) );
NOR2_X1 U16026 ( .A1(n19769), .A2(n8437), .ZN(n9300) );
NOR2_X1 U16027 ( .A1(n19757), .A2(n8150), .ZN(n8336) );
NOR2_X1 U16028 ( .A1(n19757), .A2(n8437), .ZN(n9054) );
NOR2_X1 U16029 ( .A1(n19759), .A2(n8150), .ZN(n8340) );
NOR2_X1 U16030 ( .A1(n19759), .A2(n8437), .ZN(n9095) );
NOR2_X1 U16031 ( .A1(n19761), .A2(n8150), .ZN(n8344) );
NOR2_X1 U16032 ( .A1(n19761), .A2(n8437), .ZN(n9136) );
NOR2_X1 U16033 ( .A1(n19763), .A2(n16381), .ZN(n8348) );
NOR2_X1 U16034 ( .A1(n19763), .A2(n8437), .ZN(n9177) );
NOR2_X1 U16035 ( .A1(n19765), .A2(n8150), .ZN(n8352) );
NOR2_X1 U16036 ( .A1(n19765), .A2(n8437), .ZN(n9218) );
NOR2_X1 U16037 ( .A1(n19767), .A2(n16381), .ZN(n8356) );
NOR2_X1 U16038 ( .A1(n19767), .A2(n16378), .ZN(n9259) );
NOR2_X1 U16039 ( .A1(n19771), .A2(n8150), .ZN(n8364) );
NOR2_X1 U16040 ( .A1(n19771), .A2(n8437), .ZN(n9343) );
NOR2_X1 U16041 ( .A1(n19773), .A2(n16381), .ZN(n8372) );
NOR2_X1 U16042 ( .A1(n19773), .A2(n8437), .ZN(n9430) );
NOR2_X1 U16043 ( .A1(n19775), .A2(n8150), .ZN(n8376) );
NOR2_X1 U16044 ( .A1(n19775), .A2(n16378), .ZN(n9471) );
NOR2_X1 U16045 ( .A1(n19779), .A2(n16381), .ZN(n8384) );
NOR2_X1 U16046 ( .A1(n19779), .A2(n8437), .ZN(n9556) );
NOR2_X1 U16047 ( .A1(n19781), .A2(n8150), .ZN(n8388) );
NOR2_X1 U16048 ( .A1(n19781), .A2(n16378), .ZN(n9598) );
NOR2_X1 U16049 ( .A1(n19783), .A2(n16381), .ZN(n8392) );
NOR2_X1 U16050 ( .A1(n19783), .A2(n8437), .ZN(n9636) );
NOR2_X1 U16051 ( .A1(n19785), .A2(n8150), .ZN(n8396) );
NOR2_X1 U16052 ( .A1(n19785), .A2(n16378), .ZN(n9673) );
NOR2_X1 U16053 ( .A1(n19787), .A2(n16381), .ZN(n8400) );
NOR2_X1 U16054 ( .A1(n19787), .A2(n8437), .ZN(n9710) );
NOR2_X1 U16055 ( .A1(n19789), .A2(n8150), .ZN(n8404) );
NOR2_X1 U16056 ( .A1(n19789), .A2(n16378), .ZN(n9750) );
NOR2_X1 U16057 ( .A1(n19791), .A2(n16381), .ZN(n8408) );
NOR2_X1 U16058 ( .A1(n19791), .A2(n8437), .ZN(n9798) );
NOR2_X1 U16059 ( .A1(n19807), .A2(n16378), .ZN(n8968) );
NOR2_X1 U16060 ( .A1(n19811), .A2(n16378), .ZN(n9835) );
NOR2_X1 U16061 ( .A1(n19777), .A2(n8150), .ZN(n8380) );
NOR2_X1 U16062 ( .A1(n19777), .A2(n8437), .ZN(n9512) );
NOR2_X1 U16063 ( .A1(n19755), .A2(n16381), .ZN(n8332) );
NOR2_X1 U16064 ( .A1(n19755), .A2(n8437), .ZN(n9013) );
NOR2_X1 U16065 ( .A1(n19753), .A2(n16378), .ZN(n8972) );
NOR2_X1 U16066 ( .A1(n20172), .A2(n16413), .ZN(n5421) );
NOR2_X1 U16067 ( .A1(n20749), .A2(n16413), .ZN(n5426) );
NOR2_X1 U16068 ( .A1(n20210), .A2(n16413), .ZN(n5431) );
NOR2_X1 U16069 ( .A1(n20248), .A2(n16413), .ZN(n5436) );
NOR2_X1 U16070 ( .A1(n20287), .A2(n16413), .ZN(n5440) );
NOR2_X1 U16071 ( .A1(n20326), .A2(n16413), .ZN(n5444) );
NOR2_X1 U16072 ( .A1(n20365), .A2(n16413), .ZN(n5449) );
NOR2_X1 U16073 ( .A1(n20404), .A2(n16413), .ZN(n5453) );
NOR2_X1 U16074 ( .A1(n20443), .A2(n16413), .ZN(n5457) );
NOR2_X1 U16075 ( .A1(n20483), .A2(n16413), .ZN(n5461) );
NOR2_X1 U16076 ( .A1(n20523), .A2(n16413), .ZN(n5465) );
NOR2_X1 U16077 ( .A1(n20563), .A2(n16413), .ZN(n5469) );
NOR2_X1 U16078 ( .A1(n20603), .A2(n5386), .ZN(n5478) );
NOR2_X1 U16079 ( .A1(n20641), .A2(n5386), .ZN(n5483) );
NOR2_X1 U16080 ( .A1(n20676), .A2(n5386), .ZN(n5488) );
NOR2_X1 U16081 ( .A1(n20684), .A2(n16413), .ZN(n5493) );
NOR2_X1 U16082 ( .A1(n20688), .A2(n5386), .ZN(n5498) );
NOR2_X1 U16083 ( .A1(n20692), .A2(n16413), .ZN(n5503) );
NOR2_X1 U16084 ( .A1(n20696), .A2(n5386), .ZN(n5507) );
NOR2_X1 U16085 ( .A1(n20700), .A2(n16413), .ZN(n5511) );
NOR2_X1 U16086 ( .A1(n20704), .A2(n5386), .ZN(n5516) );
NOR2_X1 U16087 ( .A1(n20708), .A2(n16413), .ZN(n5521) );
NOR2_X1 U16088 ( .A1(n20757), .A2(n5386), .ZN(n5526) );
NOR2_X1 U16089 ( .A1(n19769), .A2(n8169), .ZN(n8212) );
NOR2_X1 U16090 ( .A1(n19801), .A2(n16380), .ZN(n8284) );
NOR2_X1 U16091 ( .A1(n19807), .A2(n16380), .ZN(n8296) );
NOR2_X1 U16092 ( .A1(n19811), .A2(n16380), .ZN(n8304) );
NOR2_X1 U16093 ( .A1(n19769), .A2(n8456), .ZN(n8499) );
NOR2_X1 U16094 ( .A1(n19801), .A2(n8456), .ZN(n8732) );
NOR2_X1 U16095 ( .A1(n19807), .A2(n16377), .ZN(n8873) );
NOR2_X1 U16096 ( .A1(n19811), .A2(n8456), .ZN(n8881) );
NOR2_X1 U16097 ( .A1(n19771), .A2(n8169), .ZN(n8216) );
NOR2_X1 U16098 ( .A1(n19771), .A2(n8456), .ZN(n8503) );
NOR2_X1 U16099 ( .A1(n19773), .A2(n8169), .ZN(n8220) );
NOR2_X1 U16100 ( .A1(n19773), .A2(n8456), .ZN(n8507) );
NOR2_X1 U16101 ( .A1(n19775), .A2(n8169), .ZN(n8224) );
NOR2_X1 U16102 ( .A1(n19775), .A2(n8456), .ZN(n8511) );
NOR2_X1 U16103 ( .A1(n19779), .A2(n16380), .ZN(n8236) );
NOR2_X1 U16104 ( .A1(n19779), .A2(n8456), .ZN(n8523) );
NOR2_X1 U16105 ( .A1(n19777), .A2(n8169), .ZN(n8232) );
NOR2_X1 U16106 ( .A1(n19777), .A2(n8456), .ZN(n8519) );
NOR2_X1 U16107 ( .A1(n19765), .A2(n16380), .ZN(n8204) );
NOR2_X1 U16108 ( .A1(n19765), .A2(n8456), .ZN(n8491) );
NOR2_X1 U16109 ( .A1(n19767), .A2(n8169), .ZN(n8208) );
NOR2_X1 U16110 ( .A1(n19767), .A2(n16377), .ZN(n8495) );
NOR2_X1 U16111 ( .A1(n19781), .A2(n16380), .ZN(n8240) );
NOR2_X1 U16112 ( .A1(n19781), .A2(n8456), .ZN(n8527) );
NOR2_X1 U16113 ( .A1(n19783), .A2(n8169), .ZN(n8244) );
NOR2_X1 U16114 ( .A1(n19783), .A2(n16377), .ZN(n8531) );
NOR2_X1 U16115 ( .A1(n19785), .A2(n16380), .ZN(n8248) );
NOR2_X1 U16116 ( .A1(n19785), .A2(n8456), .ZN(n8535) );
NOR2_X1 U16117 ( .A1(n19787), .A2(n8169), .ZN(n8252) );
NOR2_X1 U16118 ( .A1(n19787), .A2(n16377), .ZN(n8539) );
NOR2_X1 U16119 ( .A1(n19789), .A2(n16380), .ZN(n8256) );
NOR2_X1 U16120 ( .A1(n19789), .A2(n16377), .ZN(n8543) );
NOR2_X1 U16121 ( .A1(n19791), .A2(n16380), .ZN(n8260) );
NOR2_X1 U16122 ( .A1(n19791), .A2(n8456), .ZN(n8547) );
NOR2_X1 U16123 ( .A1(n19793), .A2(n16380), .ZN(n8264) );
NOR2_X1 U16124 ( .A1(n19793), .A2(n16377), .ZN(n8551) );
NOR2_X1 U16125 ( .A1(n19795), .A2(n16380), .ZN(n8268) );
NOR2_X1 U16126 ( .A1(n19795), .A2(n8456), .ZN(n8604) );
NOR2_X1 U16127 ( .A1(n19799), .A2(n16380), .ZN(n8280) );
NOR2_X1 U16128 ( .A1(n19799), .A2(n16377), .ZN(n8695) );
NOR2_X1 U16129 ( .A1(n19797), .A2(n16380), .ZN(n8276) );
NOR2_X1 U16130 ( .A1(n19797), .A2(n8456), .ZN(n8647) );
NOR2_X1 U16131 ( .A1(n16440), .A2(n19823), .ZN(n3456) );
NOR2_X1 U16132 ( .A1(n16441), .A2(n19828), .ZN(n3466) );
NOR2_X1 U16133 ( .A1(n16440), .A2(n19841), .ZN(n3491) );
NOR2_X1 U16134 ( .A1(n16441), .A2(n19851), .ZN(n3522) );
NAND2_X1 U16135 ( .A1(n10505), .A2(n20964), .ZN(n6190) );
NOR2_X1 U16136 ( .A1(n4411), .A2(n4412), .ZN(n4408) );
NOR2_X1 U16137 ( .A1(n16441), .A2(n19821), .ZN(n3451) );
NAND2_X1 U16138 ( .A1(n8129), .A2(n9969), .ZN(n9891) );
NOR2_X1 U16139 ( .A1(n9925), .A2(n9908), .ZN(n9969) );
NOR2_X1 U16140 ( .A1(n19801), .A2(n16390), .ZN(n7898) );
NOR2_X1 U16141 ( .A1(n19749), .A2(n16390), .ZN(n7916) );
NOR2_X1 U16142 ( .A1(n19751), .A2(n16390), .ZN(n7922) );
NOR2_X1 U16143 ( .A1(n19769), .A2(n16391), .ZN(n7982) );
NOR2_X1 U16144 ( .A1(n19809), .A2(n16391), .ZN(n7994) );
NOR2_X1 U16145 ( .A1(n19757), .A2(n16391), .ZN(n7946) );
NOR2_X1 U16146 ( .A1(n19759), .A2(n16391), .ZN(n7952) );
NOR2_X1 U16147 ( .A1(n19761), .A2(n16391), .ZN(n7958) );
NOR2_X1 U16148 ( .A1(n19763), .A2(n16391), .ZN(n7964) );
NOR2_X1 U16149 ( .A1(n19765), .A2(n16391), .ZN(n7970) );
NOR2_X1 U16150 ( .A1(n19767), .A2(n16391), .ZN(n7976) );
NOR2_X1 U16151 ( .A1(n19771), .A2(n16391), .ZN(n7988) );
NOR2_X1 U16152 ( .A1(n19773), .A2(n16391), .ZN(n8000) );
NOR2_X1 U16153 ( .A1(n19775), .A2(n16391), .ZN(n8006) );
NOR2_X1 U16154 ( .A1(n19793), .A2(n16390), .ZN(n7870) );
NOR2_X1 U16155 ( .A1(n19795), .A2(n16390), .ZN(n7880) );
NOR2_X1 U16156 ( .A1(n19799), .A2(n16390), .ZN(n7892) );
NOR2_X1 U16157 ( .A1(n19803), .A2(n16390), .ZN(n7904) );
NOR2_X1 U16158 ( .A1(n19797), .A2(n16390), .ZN(n7886) );
NOR2_X1 U16159 ( .A1(n19805), .A2(n16390), .ZN(n7910) );
NOR2_X1 U16160 ( .A1(n19807), .A2(n16390), .ZN(n7928) );
NOR2_X1 U16161 ( .A1(n19777), .A2(n16391), .ZN(n8012) );
NOR2_X1 U16162 ( .A1(n19755), .A2(n16390), .ZN(n7940) );
NOR2_X1 U16163 ( .A1(n19753), .A2(n16390), .ZN(n7934) );
AND2_X1 U16164 ( .A1(n2343), .A2(n2344), .ZN(n2307) );
NAND2_X1 U16165 ( .A1(n16451), .A2(n2345), .ZN(n2344) );
NAND2_X1 U16166 ( .A1(n2142), .A2(n2354), .ZN(n2343) );
NAND2_X1 U16167 ( .A1(n2279), .A2(n2346), .ZN(n2345) );
NOR2_X1 U16168 ( .A1(n19797), .A2(n7052), .ZN(n7050) );
INV_X1 U16169 ( .A(n2408), .ZN(n19899) );
INV_X1 U16170 ( .A(n2222), .ZN(n19877) );
NOR2_X1 U16171 ( .A1(n2470), .A2(n2523), .ZN(n2520) );
NOR2_X1 U16172 ( .A1(n2029), .A2(n2030), .ZN(n2027) );
NOR2_X1 U16173 ( .A1(n2238), .A2(n2674), .ZN(n2673) );
NAND2_X1 U16174 ( .A1(n19888), .A2(n2557), .ZN(n2674) );
NOR2_X1 U16175 ( .A1(n19906), .A2(n19941), .ZN(n2400) );
NOR2_X1 U16176 ( .A1(n6309), .A2(n10117), .ZN(n10111) );
BUF_X1 U16177 ( .A(n3611), .Z(n16429) );
INV_X1 U16178 ( .A(n2590), .ZN(n19895) );
BUF_X1 U16179 ( .A(n3018), .Z(n16442) );
NAND2_X1 U16180 ( .A1(n2036), .A2(n2581), .ZN(n2544) );
OR2_X1 U16181 ( .A1(n2582), .A2(n16454), .ZN(n2581) );
NOR2_X1 U16182 ( .A1(n20985), .A2(n5138), .ZN(n5137) );
NAND2_X1 U16183 ( .A1(n19894), .A2(n2666), .ZN(n2141) );
NAND2_X1 U16184 ( .A1(n2236), .A2(n2237), .ZN(n2180) );
NAND2_X1 U16185 ( .A1(n2142), .A2(n2238), .ZN(n2236) );
NAND2_X1 U16186 ( .A1(n16451), .A2(n2377), .ZN(n2376) );
NAND2_X1 U16187 ( .A1(n2378), .A2(n19903), .ZN(n2377) );
NOR2_X1 U16188 ( .A1(n19889), .A2(n2026), .ZN(n2378) );
AND2_X1 U16189 ( .A1(n20945), .A2(n1394), .ZN(n1342) );
NAND2_X1 U16190 ( .A1(n20952), .A2(n6235), .ZN(n10108) );
NAND2_X1 U16191 ( .A1(n10060), .A2(n10504), .ZN(n10481) );
NOR2_X1 U16192 ( .A1(n2397), .A2(n2363), .ZN(n2768) );
NOR2_X1 U16193 ( .A1(n16455), .A2(n2113), .ZN(n2111) );
INV_X1 U16194 ( .A(n2147), .ZN(n19889) );
NAND2_X1 U16195 ( .A1(n2266), .A2(n2222), .ZN(n2265) );
INV_X1 U16196 ( .A(n2178), .ZN(n19879) );
AND2_X1 U16197 ( .A1(n7032), .A2(n20859), .ZN(n7178) );
NAND2_X1 U16198 ( .A1(n6309), .A2(n20940), .ZN(n1338) );
NAND2_X1 U16199 ( .A1(n10499), .A2(n20964), .ZN(n6186) );
NOR2_X1 U16200 ( .A1(n20966), .A2(n20956), .ZN(n10499) );
NAND2_X1 U16201 ( .A1(n8101), .A2(n16385), .ZN(n8100) );
NAND2_X1 U16202 ( .A1(n1397), .A2(n20943), .ZN(n1317) );
NOR2_X1 U16203 ( .A1(n20952), .A2(n20942), .ZN(n1397) );
NAND2_X1 U16204 ( .A1(n5225), .A2(n5143), .ZN(n3704) );
NAND2_X1 U16205 ( .A1(n2486), .A2(n19916), .ZN(n2241) );
AND2_X1 U16206 ( .A1(n2049), .A2(n2047), .ZN(n2486) );
NAND2_X1 U16207 ( .A1(n2276), .A2(n2277), .ZN(n2261) );
OR2_X1 U16208 ( .A1(n2279), .A2(n16456), .ZN(n2276) );
NAND2_X1 U16209 ( .A1(n19897), .A2(n2142), .ZN(n2277) );
AND2_X1 U16210 ( .A1(n19978), .A2(n8126), .ZN(n8086) );
NAND2_X1 U16211 ( .A1(n19809), .A2(n19811), .ZN(n8126) );
NAND2_X1 U16212 ( .A1(n2137), .A2(n2138), .ZN(n2107) );
NOR2_X1 U16213 ( .A1(n2139), .A2(n2140), .ZN(n2137) );
AND2_X1 U16214 ( .A1(n2141), .A2(n2142), .ZN(n2140) );
AND2_X1 U16215 ( .A1(n1401), .A2(n1394), .ZN(n1315) );
NOR2_X1 U16216 ( .A1(n20945), .A2(n20944), .ZN(n1401) );
INV_X1 U16217 ( .A(n2055), .ZN(n19902) );
AND2_X1 U16218 ( .A1(n2380), .A2(n2381), .ZN(n2009) );
NAND2_X1 U16219 ( .A1(n16451), .A2(n2382), .ZN(n2381) );
NAND2_X1 U16220 ( .A1(n2142), .A2(n2184), .ZN(n2380) );
NAND2_X1 U16221 ( .A1(n2383), .A2(n2384), .ZN(n2382) );
AND2_X1 U16222 ( .A1(n8097), .A2(n8098), .ZN(n7082) );
NOR2_X1 U16223 ( .A1(n8107), .A2(n8108), .ZN(n8097) );
NOR2_X1 U16224 ( .A1(n8099), .A2(n8100), .ZN(n8098) );
NAND2_X1 U16225 ( .A1(n20832), .A2(n20860), .ZN(n8108) );
AND2_X1 U16226 ( .A1(n2534), .A2(n2535), .ZN(n2078) );
NAND2_X1 U16227 ( .A1(n19898), .A2(n16453), .ZN(n2535) );
NOR2_X1 U16228 ( .A1(n2536), .A2(n2537), .ZN(n2534) );
NOR2_X1 U16229 ( .A1(n2352), .A2(n2457), .ZN(n2536) );
NAND2_X1 U16230 ( .A1(n1404), .A2(n20940), .ZN(n1335) );
NOR2_X1 U16231 ( .A1(n20952), .A2(n16468), .ZN(n1404) );
NAND2_X1 U16232 ( .A1(n2363), .A2(n16450), .ZN(n2360) );
INV_X1 U16233 ( .A(n10501), .ZN(n20966) );
AND2_X1 U16234 ( .A1(n2691), .A2(n2692), .ZN(n2367) );
NOR2_X1 U16235 ( .A1(n2693), .A2(n2694), .ZN(n2692) );
NOR2_X1 U16236 ( .A1(n2698), .A2(n2699), .ZN(n2691) );
NOR2_X1 U16237 ( .A1(n16457), .A2(n2695), .ZN(n2693) );
AND2_X1 U16238 ( .A1(n2474), .A2(n2475), .ZN(n2066) );
NOR2_X1 U16239 ( .A1(n2481), .A2(n2482), .ZN(n2474) );
NAND2_X1 U16240 ( .A1(n2142), .A2(n2476), .ZN(n2475) );
NOR2_X1 U16241 ( .A1(n2483), .A2(n16456), .ZN(n2481) );
AND2_X1 U16242 ( .A1(n2707), .A2(n2708), .ZN(n2370) );
NOR2_X1 U16243 ( .A1(n2721), .A2(n2722), .ZN(n2707) );
NAND2_X1 U16244 ( .A1(n2142), .A2(n2709), .ZN(n2708) );
NOR2_X1 U16245 ( .A1(n2725), .A2(n16456), .ZN(n2721) );
INV_X1 U16246 ( .A(n2557), .ZN(n19900) );
AND2_X1 U16247 ( .A1(n2682), .A2(n2142), .ZN(n2699) );
INV_X1 U16248 ( .A(n2113), .ZN(n19890) );
INV_X1 U16249 ( .A(n6235), .ZN(n20942) );
INV_X1 U16250 ( .A(n2363), .ZN(n19903) );
INV_X1 U16251 ( .A(n5143), .ZN(n20983) );
INV_X1 U16252 ( .A(n2339), .ZN(n19880) );
INV_X1 U16253 ( .A(n2453), .ZN(n19888) );
INV_X1 U16254 ( .A(n10504), .ZN(n20954) );
INV_X1 U16255 ( .A(n2048), .ZN(n19916) );
NAND2_X1 U16256 ( .A1(n8103), .A2(n16383), .ZN(n8099) );
NOR2_X1 U16257 ( .A1(n7795), .A2(n20844), .ZN(n8103) );
NAND2_X1 U16258 ( .A1(n2269), .A2(n2696), .ZN(n2695) );
AND2_X1 U16259 ( .A1(n8165), .A2(n8306), .ZN(n8168) );
INV_X1 U16260 ( .A(n2384), .ZN(n19898) );
INV_X1 U16261 ( .A(n4936), .ZN(n20909) );
NAND2_X1 U16262 ( .A1(n2355), .A2(n2356), .ZN(n2354) );
NOR2_X1 U16263 ( .A1(n19897), .A2(n19891), .ZN(n2355) );
OR2_X1 U16264 ( .A1(n20725), .A2(n21395), .ZN(n21396) );
OR2_X1 U16265 ( .A1(n19870), .A2(n21401), .ZN(n21402) );
OR2_X1 U16266 ( .A1(n19865), .A2(n21311), .ZN(n21308) );
OR2_X1 U16267 ( .A1(n19860), .A2(n21318), .ZN(n21315) );
OR2_X1 U16268 ( .A1(n19855), .A2(n21325), .ZN(n21322) );
OR2_X1 U16269 ( .A1(n19850), .A2(n21332), .ZN(n21329) );
OR2_X1 U16270 ( .A1(n19845), .A2(n21339), .ZN(n21336) );
OR2_X1 U16271 ( .A1(n19840), .A2(n21346), .ZN(n21343) );
OR2_X1 U16272 ( .A1(n19835), .A2(n21353), .ZN(n21350) );
OR2_X1 U16273 ( .A1(n19830), .A2(n21360), .ZN(n21357) );
OR2_X1 U16274 ( .A1(n19825), .A2(n21367), .ZN(n21364) );
OR2_X1 U16275 ( .A1(n19820), .A2(n21376), .ZN(n21371) );
OR2_X1 U16276 ( .A1(n20736), .A2(n21389), .ZN(n21390) );
NAND2_X1 U16277 ( .A1(n20878), .A2(n20747), .ZN(n21374) );
AND2_X1 U16278 ( .A1(n4275), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_8), .ZN(n4294) );
AND2_X1 U16279 ( .A1(n2461), .A2(n2728), .ZN(n2669) );
NAND2_X1 U16280 ( .A1(n16450), .A2(n2184), .ZN(n2728) );
AND2_X1 U16281 ( .A1(n2048), .A2(n2049), .ZN(n2046) );
INV_X1 U16282 ( .A(n8414), .ZN(n19979) );
INV_X1 U16283 ( .A(n10127), .ZN(n20941) );
INV_X1 U16284 ( .A(n4049), .ZN(n20874) );
NOR2_X1 U16285 ( .A1(n21259), .A2(n21258), .ZN(data_addr_o_31_) );
AND2_X1 U16286 ( .A1(n21257), .A2(n21256), .ZN(n21258) );
NAND2_X1 U16287 ( .A1(n21251), .A2(n21250), .ZN(n21256) );
NAND2_X1 U16288 ( .A1(n21080), .A2(n21079), .ZN(n21086) );
NAND2_X1 U16289 ( .A1(ex_block_i_alu_i_adder_in_a_13), .A2(n21077), .ZN(n21080) );
OR2_X1 U16290 ( .A1(n21077), .A2(ex_block_i_alu_i_adder_in_a_13), .ZN(n21078) );
NAND2_X1 U16291 ( .A1(n21098), .A2(n21097), .ZN(n21104) );
NAND2_X1 U16292 ( .A1(ex_block_i_alu_i_adder_in_a_15), .A2(n21095), .ZN(n21098) );
OR2_X1 U16293 ( .A1(n21095), .A2(ex_block_i_alu_i_adder_in_a_15), .ZN(n21096) );
NAND2_X1 U16294 ( .A1(n21107), .A2(n21106), .ZN(n21113) );
NAND2_X1 U16295 ( .A1(ex_block_i_alu_i_adder_in_a_16), .A2(n21104), .ZN(n21107) );
OR2_X1 U16296 ( .A1(n21104), .A2(ex_block_i_alu_i_adder_in_a_16), .ZN(n21105) );
NAND2_X1 U16297 ( .A1(n21139), .A2(n21138), .ZN(n21145) );
NAND2_X1 U16298 ( .A1(ex_block_i_alu_i_adder_in_a_19), .A2(n21136), .ZN(n21139) );
OR2_X1 U16299 ( .A1(n21136), .A2(ex_block_i_alu_i_adder_in_a_19), .ZN(n21137) );
NAND2_X1 U16300 ( .A1(n21148), .A2(n21147), .ZN(n21154) );
NAND2_X1 U16301 ( .A1(ex_block_i_alu_i_adder_in_a_20), .A2(n21145), .ZN(n21148) );
OR2_X1 U16302 ( .A1(n21145), .A2(ex_block_i_alu_i_adder_in_a_20), .ZN(n21146) );
NAND2_X1 U16303 ( .A1(n21166), .A2(n21165), .ZN(n21172) );
NAND2_X1 U16304 ( .A1(ex_block_i_alu_i_adder_in_a_22), .A2(n21163), .ZN(n21166) );
OR2_X1 U16305 ( .A1(n21163), .A2(ex_block_i_alu_i_adder_in_a_22), .ZN(n21164) );
NAND2_X1 U16306 ( .A1(n21175), .A2(n21174), .ZN(n21181) );
NAND2_X1 U16307 ( .A1(ex_block_i_alu_i_adder_in_a_23), .A2(n21172), .ZN(n21175) );
OR2_X1 U16308 ( .A1(n21172), .A2(ex_block_i_alu_i_adder_in_a_23), .ZN(n21173) );
NAND2_X1 U16309 ( .A1(n21193), .A2(n21192), .ZN(n21199) );
NAND2_X1 U16310 ( .A1(ex_block_i_alu_i_adder_in_a_25), .A2(n21190), .ZN(n21193) );
OR2_X1 U16311 ( .A1(n21190), .A2(ex_block_i_alu_i_adder_in_a_25), .ZN(n21191) );
NAND2_X1 U16312 ( .A1(n21202), .A2(n21201), .ZN(n21208) );
NAND2_X1 U16313 ( .A1(ex_block_i_alu_i_adder_in_a_26), .A2(n21199), .ZN(n21202) );
OR2_X1 U16314 ( .A1(n21199), .A2(ex_block_i_alu_i_adder_in_a_26), .ZN(n21200) );
NAND2_X1 U16315 ( .A1(n21235), .A2(n21234), .ZN(n21241) );
NAND2_X1 U16316 ( .A1(ex_block_i_alu_i_adder_in_a_29), .A2(n21232), .ZN(n21235) );
OR2_X1 U16317 ( .A1(n21232), .A2(ex_block_i_alu_i_adder_in_a_29), .ZN(n21233) );
NOR2_X1 U16318 ( .A1(n20939), .A2(n20869), .ZN(n5938) );
NOR2_X1 U16319 ( .A1(n20939), .A2(n20871), .ZN(n6090) );
NOR2_X1 U16320 ( .A1(n20939), .A2(n20864), .ZN(n5884) );
NOR2_X1 U16321 ( .A1(n20939), .A2(n20861), .ZN(n5874) );
NOR2_X1 U16322 ( .A1(n20939), .A2(n20853), .ZN(n5864) );
NAND2_X1 U16323 ( .A1(n21244), .A2(n21243), .ZN(n21252) );
NAND2_X1 U16324 ( .A1(ex_block_i_alu_i_adder_in_a_30), .A2(n21241), .ZN(n21244) );
OR2_X1 U16325 ( .A1(n21241), .A2(ex_block_i_alu_i_adder_in_a_30), .ZN(n21242) );
NAND2_X1 U16326 ( .A1(n21089), .A2(n21088), .ZN(n21095) );
NAND2_X1 U16327 ( .A1(ex_block_i_alu_i_adder_in_a_14), .A2(n21086), .ZN(n21089) );
NAND2_X1 U16328 ( .A1(ex_block_i_alu_i_adder_in_b_14), .A2(n21087), .ZN(n21088) );
OR2_X1 U16329 ( .A1(n21086), .A2(ex_block_i_alu_i_adder_in_a_14), .ZN(n21087) );
NAND2_X1 U16330 ( .A1(n21116), .A2(n21115), .ZN(n21122) );
NAND2_X1 U16331 ( .A1(ex_block_i_alu_i_adder_in_a_17), .A2(n21113), .ZN(n21116) );
NAND2_X1 U16332 ( .A1(ex_block_i_alu_i_adder_in_b_17), .A2(n21114), .ZN(n21115) );
OR2_X1 U16333 ( .A1(n21113), .A2(ex_block_i_alu_i_adder_in_a_17), .ZN(n21114) );
NAND2_X1 U16334 ( .A1(n21125), .A2(n21124), .ZN(n21136) );
NAND2_X1 U16335 ( .A1(ex_block_i_alu_i_adder_in_a_18), .A2(n21122), .ZN(n21125) );
NAND2_X1 U16336 ( .A1(ex_block_i_alu_i_adder_in_b_18), .A2(n21123), .ZN(n21124) );
OR2_X1 U16337 ( .A1(n21122), .A2(ex_block_i_alu_i_adder_in_a_18), .ZN(n21123) );
NAND2_X1 U16338 ( .A1(n21157), .A2(n21156), .ZN(n21163) );
NAND2_X1 U16339 ( .A1(ex_block_i_alu_i_adder_in_a_21), .A2(n21154), .ZN(n21157) );
NAND2_X1 U16340 ( .A1(ex_block_i_alu_i_adder_in_b_21), .A2(n21155), .ZN(n21156) );
OR2_X1 U16341 ( .A1(n21154), .A2(ex_block_i_alu_i_adder_in_a_21), .ZN(n21155) );
NAND2_X1 U16342 ( .A1(n21184), .A2(n21183), .ZN(n21190) );
NAND2_X1 U16343 ( .A1(ex_block_i_alu_i_adder_in_a_24), .A2(n21181), .ZN(n21184) );
NAND2_X1 U16344 ( .A1(ex_block_i_alu_i_adder_in_b_24), .A2(n21182), .ZN(n21183) );
OR2_X1 U16345 ( .A1(n21181), .A2(ex_block_i_alu_i_adder_in_a_24), .ZN(n21182) );
NAND2_X1 U16346 ( .A1(n21211), .A2(n21210), .ZN(n21217) );
NAND2_X1 U16347 ( .A1(ex_block_i_alu_i_adder_in_a_27), .A2(n21208), .ZN(n21211) );
NAND2_X1 U16348 ( .A1(ex_block_i_alu_i_adder_in_b_27), .A2(n21209), .ZN(n21210) );
OR2_X1 U16349 ( .A1(n21208), .A2(ex_block_i_alu_i_adder_in_a_27), .ZN(n21209) );
NAND2_X1 U16350 ( .A1(n21220), .A2(n21219), .ZN(n21232) );
NAND2_X1 U16351 ( .A1(ex_block_i_alu_i_adder_in_a_28), .A2(n21217), .ZN(n21220) );
NAND2_X1 U16352 ( .A1(ex_block_i_alu_i_adder_in_b_28), .A2(n21218), .ZN(n21219) );
OR2_X1 U16353 ( .A1(n21217), .A2(ex_block_i_alu_i_adder_in_a_28), .ZN(n21218) );
NOR2_X1 U16354 ( .A1(n20112), .A2(n10115), .ZN(n10121) );
NOR2_X1 U16355 ( .A1(n19815), .A2(n16458), .ZN(n1754) );
NOR2_X1 U16356 ( .A1(n19813), .A2(n1708), .ZN(n1748) );
AND2_X1 U16357 ( .A1(n5272), .A2(n4257), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_sign_b) );
NOR2_X1 U16358 ( .A1(n6310), .A2(n10090), .ZN(n10087) );
NAND2_X1 U16359 ( .A1(n20952), .A2(n20111), .ZN(n10090) );
NOR2_X1 U16360 ( .A1(n10119), .A2(n10120), .ZN(n10105) );
NOR2_X1 U16361 ( .A1(n6234), .A2(n10159), .ZN(n10119) );
NOR2_X1 U16362 ( .A1(n10121), .A2(n10122), .ZN(n10120) );
NAND2_X1 U16363 ( .A1(n10160), .A2(n10127), .ZN(n10159) );
NOR2_X1 U16364 ( .A1(n10113), .A2(n10114), .ZN(n10112) );
AND2_X1 U16365 ( .A1(n10115), .A2(n10116), .ZN(n10114) );
NOR2_X1 U16366 ( .A1(data_addr_o_31_), .A2(n10115), .ZN(n10113) );
NAND2_X1 U16367 ( .A1(n16471), .A2(n1415), .ZN(n1378) );
NAND2_X1 U16368 ( .A1(n20819), .A2(n1380), .ZN(n1379) );
NAND2_X1 U16369 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
INV_X1 U16370 ( .A(ex_block_i_alu_i_adder_in_a_1), .ZN(n20758) );
NAND2_X1 U16371 ( .A1(n21255), .A2(n21254), .ZN(n21257) );
NAND2_X1 U16372 ( .A1(ex_block_i_alu_i_adder_in_a_31), .A2(n21252), .ZN(n21255) );
NAND2_X1 U16373 ( .A1(ex_block_i_alu_i_adder_in_b_31), .A2(n21253), .ZN(n21254) );
OR2_X1 U16374 ( .A1(n21252), .A2(ex_block_i_alu_i_adder_in_a_31), .ZN(n21253) );
NOR2_X1 U16375 ( .A1(n20939), .A2(n20846), .ZN(n5854) );
NOR2_X1 U16376 ( .A1(n20939), .A2(n20841), .ZN(n5844) );
NOR2_X1 U16377 ( .A1(n20939), .A2(n20839), .ZN(n5833) );
NOR2_X1 U16378 ( .A1(n20939), .A2(n20835), .ZN(n5820) );
NOR2_X1 U16379 ( .A1(n20939), .A2(n20833), .ZN(n6223) );
NOR2_X1 U16380 ( .A1(n20939), .A2(n20830), .ZN(n6211) );
NOR2_X1 U16381 ( .A1(n19831), .A2(n16458), .ZN(n1796) );
NOR2_X1 U16382 ( .A1(n19828), .A2(n16458), .ZN(n1790) );
NOR2_X1 U16383 ( .A1(n19826), .A2(n16458), .ZN(n1784) );
NOR2_X1 U16384 ( .A1(n19823), .A2(n16458), .ZN(n1778) );
NOR2_X1 U16385 ( .A1(n19821), .A2(n1708), .ZN(n1772) );
NOR2_X1 U16386 ( .A1(n19818), .A2(n1708), .ZN(n1766) );
INV_X1 U16387 ( .A(n3467), .ZN(n19828) );
INV_X1 U16388 ( .A(n3457), .ZN(n19823) );
INV_X1 U16389 ( .A(n3452), .ZN(n19821) );
NOR2_X1 U16390 ( .A1(n20939), .A2(n20828), .ZN(n6201) );
NOR2_X1 U16391 ( .A1(n19846), .A2(n16458), .ZN(n1832) );
NOR2_X1 U16392 ( .A1(n19843), .A2(n16458), .ZN(n1826) );
NOR2_X1 U16393 ( .A1(n19841), .A2(n16458), .ZN(n1820) );
NOR2_X1 U16394 ( .A1(n19838), .A2(n16458), .ZN(n1814) );
NOR2_X1 U16395 ( .A1(n19836), .A2(n16458), .ZN(n1808) );
NOR2_X1 U16396 ( .A1(n19833), .A2(n16458), .ZN(n1802) );
INV_X1 U16397 ( .A(n3492), .ZN(n19841) );
NAND2_X1 U16398 ( .A1(n1200), .A2(n1201), .ZN(n1193) );
NAND2_X1 U16399 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_18), .A2(n87), .ZN(n1201) );
NOR2_X1 U16400 ( .A1(n1202), .A2(n1203), .ZN(n1200) );
NOR2_X1 U16401 ( .A1(n90), .A2(n20696), .ZN(n1203) );
NAND2_X1 U16402 ( .A1(n1161), .A2(n1162), .ZN(n1154) );
NAND2_X1 U16403 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_17), .A2(n87), .ZN(n1162) );
NOR2_X1 U16404 ( .A1(n1163), .A2(n1164), .ZN(n1161) );
NOR2_X1 U16405 ( .A1(n90), .A2(n20692), .ZN(n1164) );
NAND2_X1 U16406 ( .A1(n1122), .A2(n1123), .ZN(n1115) );
NAND2_X1 U16407 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_16), .A2(n87), .ZN(n1123) );
NOR2_X1 U16408 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
NOR2_X1 U16409 ( .A1(n90), .A2(n20688), .ZN(n1125) );
NOR2_X1 U16410 ( .A1(n21067), .A2(n21066), .ZN(data_addr_o_11_) );
AND2_X1 U16411 ( .A1(n21068), .A2(n21065), .ZN(n21066) );
NOR2_X1 U16412 ( .A1(n21068), .A2(n21065), .ZN(n21067) );
NAND2_X1 U16413 ( .A1(n21064), .A2(n21063), .ZN(n21065) );
NOR2_X1 U16414 ( .A1(n21049), .A2(n21048), .ZN(data_addr_o_9_) );
NOR2_X1 U16415 ( .A1(n21050), .A2(n21047), .ZN(n21049) );
AND2_X1 U16416 ( .A1(n21050), .A2(n21047), .ZN(n21048) );
NAND2_X1 U16417 ( .A1(n21046), .A2(n21045), .ZN(n21047) );
NOR2_X1 U16418 ( .A1(n21058), .A2(n21057), .ZN(data_addr_o_10_) );
NOR2_X1 U16419 ( .A1(n21059), .A2(n21056), .ZN(n21058) );
AND2_X1 U16420 ( .A1(n21059), .A2(n21056), .ZN(n21057) );
NAND2_X1 U16421 ( .A1(n21055), .A2(n21054), .ZN(n21056) );
NOR2_X1 U16422 ( .A1(n21076), .A2(n21075), .ZN(data_addr_o_12_) );
NOR2_X1 U16423 ( .A1(n21077), .A2(n21074), .ZN(n21076) );
AND2_X1 U16424 ( .A1(n21077), .A2(n21074), .ZN(n21075) );
NAND2_X1 U16425 ( .A1(n21073), .A2(n21072), .ZN(n21074) );
NOR2_X1 U16426 ( .A1(n19861), .A2(n16458), .ZN(n1868) );
NOR2_X1 U16427 ( .A1(n19858), .A2(n1708), .ZN(n1862) );
NOR2_X1 U16428 ( .A1(n19856), .A2(n1708), .ZN(n1856) );
NOR2_X1 U16429 ( .A1(n19853), .A2(n1708), .ZN(n1850) );
NOR2_X1 U16430 ( .A1(n19851), .A2(n16458), .ZN(n1844) );
NOR2_X1 U16431 ( .A1(n19848), .A2(n16458), .ZN(n1838) );
INV_X1 U16432 ( .A(n3523), .ZN(n19851) );
AND2_X1 U16433 ( .A1(n5274), .A2(n20085), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_sign_a) );
NAND2_X1 U16434 ( .A1(n85), .A2(n86), .ZN(n74) );
NAND2_X1 U16435 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_22), .A2(n87), .ZN(n86) );
NOR2_X1 U16436 ( .A1(n88), .A2(n89), .ZN(n85) );
NOR2_X1 U16437 ( .A1(n16469), .A2(n20712), .ZN(n89) );
NAND2_X1 U16438 ( .A1(n1336), .A2(n1337), .ZN(n1327) );
NAND2_X1 U16439 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_21), .A2(n87), .ZN(n1337) );
NOR2_X1 U16440 ( .A1(n1339), .A2(n1340), .ZN(n1336) );
NOR2_X1 U16441 ( .A1(n90), .A2(n20708), .ZN(n1340) );
NAND2_X1 U16442 ( .A1(n1278), .A2(n1279), .ZN(n1271) );
NAND2_X1 U16443 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_20), .A2(n87), .ZN(n1279) );
NOR2_X1 U16444 ( .A1(n1280), .A2(n1281), .ZN(n1278) );
NOR2_X1 U16445 ( .A1(n90), .A2(n20704), .ZN(n1281) );
NAND2_X1 U16446 ( .A1(n1239), .A2(n1240), .ZN(n1232) );
NAND2_X1 U16447 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_19), .A2(n87), .ZN(n1240) );
NOR2_X1 U16448 ( .A1(n1241), .A2(n1242), .ZN(n1239) );
NOR2_X1 U16449 ( .A1(n90), .A2(n20700), .ZN(n1242) );
NAND2_X1 U16450 ( .A1(n1413), .A2(n20962), .ZN(n386) );
NAND2_X1 U16451 ( .A1(n1422), .A2(n1419), .ZN(n359) );
NAND2_X1 U16452 ( .A1(n1419), .A2(n1420), .ZN(n92) );
NOR2_X1 U16453 ( .A1(n21271), .A2(n21270), .ZN(data_addr_o_3_) );
NOR2_X1 U16454 ( .A1(n21269), .A2(n21268), .ZN(n21271) );
AND2_X1 U16455 ( .A1(n21269), .A2(n21268), .ZN(n21270) );
NAND2_X1 U16456 ( .A1(n21267), .A2(n21266), .ZN(n21268) );
NOR2_X1 U16457 ( .A1(n21283), .A2(n21282), .ZN(data_addr_o_5_) );
NOR2_X1 U16458 ( .A1(n21281), .A2(n21280), .ZN(n21283) );
AND2_X1 U16459 ( .A1(n21281), .A2(n21280), .ZN(n21282) );
NAND2_X1 U16460 ( .A1(n21279), .A2(n21278), .ZN(n21280) );
NOR2_X1 U16461 ( .A1(n21295), .A2(n21294), .ZN(data_addr_o_7_) );
NOR2_X1 U16462 ( .A1(n21293), .A2(n21292), .ZN(n21295) );
AND2_X1 U16463 ( .A1(n21293), .A2(n21292), .ZN(n21294) );
NAND2_X1 U16464 ( .A1(n21291), .A2(n21290), .ZN(n21292) );
NOR2_X1 U16465 ( .A1(n21277), .A2(n21276), .ZN(data_addr_o_4_) );
NOR2_X1 U16466 ( .A1(n21275), .A2(n21274), .ZN(n21277) );
AND2_X1 U16467 ( .A1(n21275), .A2(n21274), .ZN(n21276) );
NAND2_X1 U16468 ( .A1(n21273), .A2(n21272), .ZN(n21274) );
NOR2_X1 U16469 ( .A1(n21289), .A2(n21288), .ZN(data_addr_o_6_) );
NOR2_X1 U16470 ( .A1(n21287), .A2(n21286), .ZN(n21289) );
AND2_X1 U16471 ( .A1(n21287), .A2(n21286), .ZN(n21288) );
NAND2_X1 U16472 ( .A1(n21285), .A2(n21284), .ZN(n21286) );
NOR2_X1 U16473 ( .A1(n21301), .A2(n21300), .ZN(data_addr_o_8_) );
NOR2_X1 U16474 ( .A1(n21299), .A2(n21298), .ZN(n21301) );
AND2_X1 U16475 ( .A1(n21299), .A2(n21298), .ZN(n21300) );
NAND2_X1 U16476 ( .A1(n21297), .A2(n21296), .ZN(n21298) );
NOR2_X1 U16477 ( .A1(n20871), .A2(n20869), .ZN(n7033) );
NAND2_X1 U16478 ( .A1(n20864), .A2(n20861), .ZN(n9918) );
NOR2_X1 U16479 ( .A1(n20937), .A2(n32), .ZN(n1413) );
INV_X1 U16480 ( .A(n10043), .ZN(n20845) );
INV_X1 U16481 ( .A(n9970), .ZN(n20838) );
NAND2_X1 U16482 ( .A1(n20838), .A2(n20841), .ZN(n9841) );
NOR2_X1 U16483 ( .A1(n16250), .A2(n16251), .ZN(n9984) );
NAND2_X1 U16484 ( .A1(n20845), .A2(n8106), .ZN(n16250) );
OR2_X1 U16485 ( .A1(n20853), .A2(n9918), .ZN(n16251) );
NOR2_X1 U16486 ( .A1(n15795), .A2(n286), .ZN(n283) );
NOR2_X1 U16487 ( .A1(n20853), .A2(n15794), .ZN(n286) );
NOR2_X1 U16488 ( .A1(n19866), .A2(n1708), .ZN(n1880) );
NOR2_X1 U16489 ( .A1(n19863), .A2(n1708), .ZN(n1874) );
NOR2_X1 U16490 ( .A1(n20726), .A2(n1708), .ZN(n1724) );
NOR2_X1 U16491 ( .A1(n20720), .A2(n1708), .ZN(n1718) );
NOR2_X1 U16492 ( .A1(n19871), .A2(n1708), .ZN(n1712) );
NOR2_X1 U16493 ( .A1(n19868), .A2(n1708), .ZN(n1704) );
NAND2_X1 U16494 ( .A1(n7719), .A2(n9984), .ZN(n8102) );
NAND2_X1 U16495 ( .A1(n20871), .A2(n20869), .ZN(n9927) );
INV_X1 U16496 ( .A(n3548), .ZN(n19863) );
NOR2_X1 U16497 ( .A1(n8106), .A2(n9998), .ZN(n9996) );
NOR2_X1 U16498 ( .A1(n9918), .A2(n9999), .ZN(n9998) );
NAND2_X1 U16499 ( .A1(n10000), .A2(n9970), .ZN(n9999) );
OR2_X1 U16500 ( .A1(n7571), .A2(n7719), .ZN(n10000) );
NOR2_X1 U16501 ( .A1(n15795), .A2(n887), .ZN(n884) );
NOR2_X1 U16502 ( .A1(n20869), .A2(n15794), .ZN(n887) );
NOR2_X1 U16503 ( .A1(n15795), .A2(n327), .ZN(n324) );
NOR2_X1 U16504 ( .A1(n20861), .A2(n15794), .ZN(n327) );
NAND2_X1 U16505 ( .A1(n16475), .A2(n20869), .ZN(n885) );
NAND2_X1 U16506 ( .A1(n20827), .A2(n7571), .ZN(n10008) );
NAND2_X1 U16507 ( .A1(n9984), .A2(n7571), .ZN(n8104) );
INV_X1 U16508 ( .A(n7581), .ZN(n20881) );
NAND2_X1 U16509 ( .A1(n16475), .A2(n20861), .ZN(n325) );
NAND2_X1 U16510 ( .A1(n16474), .A2(n20853), .ZN(n284) );
INV_X1 U16511 ( .A(n8430), .ZN(n20822) );
NAND2_X1 U16512 ( .A1(n264), .A2(n265), .ZN(n256) );
NAND2_X1 U16513 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_26), .A2(n87), .ZN(n265) );
NOR2_X1 U16514 ( .A1(n266), .A2(n267), .ZN(n264) );
NOR2_X1 U16515 ( .A1(n16469), .A2(n20732), .ZN(n267) );
NAND2_X1 U16516 ( .A1(n222), .A2(n223), .ZN(n214) );
NAND2_X1 U16517 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_25), .A2(n87), .ZN(n223) );
NOR2_X1 U16518 ( .A1(n224), .A2(n225), .ZN(n222) );
NOR2_X1 U16519 ( .A1(n16469), .A2(n20727), .ZN(n225) );
NAND2_X1 U16520 ( .A1(n179), .A2(n180), .ZN(n171) );
NAND2_X1 U16521 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_24), .A2(n87), .ZN(n180) );
NOR2_X1 U16522 ( .A1(n181), .A2(n182), .ZN(n179) );
NOR2_X1 U16523 ( .A1(n16469), .A2(n20721), .ZN(n182) );
NAND2_X1 U16524 ( .A1(n131), .A2(n132), .ZN(n123) );
NAND2_X1 U16525 ( .A1(ex_block_i_alu_i_shift_result_ext_signed_23), .A2(n87), .ZN(n132) );
NOR2_X1 U16526 ( .A1(n133), .A2(n134), .ZN(n131) );
NOR2_X1 U16527 ( .A1(n16469), .A2(n20716), .ZN(n134) );
NAND2_X1 U16528 ( .A1(n20880), .A2(n5164), .ZN(n10322) );
NAND2_X1 U16529 ( .A1(n880), .A2(n881), .ZN(n873) );
NAND2_X1 U16530 ( .A1(n882), .A2(n883), .ZN(n881) );
NOR2_X1 U16531 ( .A1(n888), .A2(n889), .ZN(n880) );
NAND2_X1 U16532 ( .A1(n884), .A2(n885), .ZN(n882) );
NAND2_X1 U16533 ( .A1(n320), .A2(n321), .ZN(n313) );
NAND2_X1 U16534 ( .A1(n322), .A2(n323), .ZN(n321) );
NOR2_X1 U16535 ( .A1(n328), .A2(n329), .ZN(n320) );
NAND2_X1 U16536 ( .A1(n324), .A2(n325), .ZN(n322) );
NAND2_X1 U16537 ( .A1(n279), .A2(n280), .ZN(n272) );
NAND2_X1 U16538 ( .A1(n281), .A2(n282), .ZN(n280) );
NOR2_X1 U16539 ( .A1(n287), .A2(n288), .ZN(n279) );
NAND2_X1 U16540 ( .A1(n283), .A2(n284), .ZN(n281) );
NAND2_X1 U16541 ( .A1(n9993), .A2(n9994), .ZN(n9977) );
NAND2_X1 U16542 ( .A1(n20844), .A2(n9995), .ZN(n9994) );
NOR2_X1 U16543 ( .A1(n10003), .A2(n10004), .ZN(n9993) );
NAND2_X1 U16544 ( .A1(n9996), .A2(n9997), .ZN(n9995) );
NAND2_X1 U16545 ( .A1(n452), .A2(n453), .ZN(n451) );
NOR2_X1 U16546 ( .A1(n15795), .A2(n455), .ZN(n452) );
NAND2_X1 U16547 ( .A1(n20751), .A2(n16474), .ZN(n453) );
NOR2_X1 U16548 ( .A1(n20751), .A2(n15794), .ZN(n455) );
NAND2_X1 U16549 ( .A1(n241), .A2(n242), .ZN(n239) );
NOR2_X1 U16550 ( .A1(n15795), .A2(n244), .ZN(n241) );
NAND2_X1 U16551 ( .A1(n20846), .A2(n16474), .ZN(n242) );
NOR2_X1 U16552 ( .A1(n20846), .A2(n15794), .ZN(n244) );
NAND2_X1 U16553 ( .A1(n198), .A2(n199), .ZN(n196) );
NOR2_X1 U16554 ( .A1(n15795), .A2(n201), .ZN(n198) );
NAND2_X1 U16555 ( .A1(n20729), .A2(n16474), .ZN(n199) );
NOR2_X1 U16556 ( .A1(n20729), .A2(n15794), .ZN(n201) );
NAND2_X1 U16557 ( .A1(n150), .A2(n151), .ZN(n148) );
NOR2_X1 U16558 ( .A1(n15795), .A2(n154), .ZN(n150) );
NAND2_X1 U16559 ( .A1(n20723), .A2(n16474), .ZN(n151) );
NOR2_X1 U16560 ( .A1(n20723), .A2(n15794), .ZN(n154) );
NOR2_X1 U16561 ( .A1(n21265), .A2(n21264), .ZN(data_addr_o_2_) );
NOR2_X1 U16562 ( .A1(n21263), .A2(n21262), .ZN(n21265) );
AND2_X1 U16563 ( .A1(n21263), .A2(n21262), .ZN(n21264) );
NAND2_X1 U16564 ( .A1(n21261), .A2(n21260), .ZN(n21262) );
INV_X1 U16565 ( .A(n10002), .ZN(n20827) );
NAND2_X1 U16566 ( .A1(ex_block_i_alu_i_shift_amt_3), .A2(n20863), .ZN(n21949) );
NOR2_X1 U16567 ( .A1(n9782), .A2(n20843), .ZN(n9938) );
NAND2_X1 U16568 ( .A1(n9938), .A2(n7719), .ZN(n8806) );
NAND2_X1 U16569 ( .A1(n10043), .A2(n20853), .ZN(n8121) );
NOR2_X1 U16570 ( .A1(ex_block_i_alu_i_shift_amt_0), .A2(ex_block_i_alu_i_shift_amt_1), .ZN(n21773) );
NAND2_X1 U16571 ( .A1(n20838), .A2(n10002), .ZN(n8115) );
NAND2_X1 U16572 ( .A1(n9780), .A2(n20858), .ZN(n8677) );
NOR2_X1 U16573 ( .A1(n8121), .A2(n9782), .ZN(n9780) );
NAND2_X1 U16574 ( .A1(ex_block_i_alu_i_shift_amt_2), .A2(n21706), .ZN(n22009) );
NOR2_X1 U16575 ( .A1(n7613), .A2(n20881), .ZN(n4036) );
AND2_X1 U16576 ( .A1(n7615), .A2(n7616), .ZN(n7613) );
NOR2_X1 U16577 ( .A1(n7617), .A2(n7618), .ZN(n7616) );
NOR2_X1 U16578 ( .A1(n20886), .A2(n7625), .ZN(n7615) );
NOR2_X1 U16579 ( .A1(n8121), .A2(n9924), .ZN(n9789) );
NAND2_X1 U16580 ( .A1(n20841), .A2(n9970), .ZN(n9908) );
NOR2_X1 U16581 ( .A1(n20856), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n21706) );
NAND2_X1 U16582 ( .A1(ex_block_i_alu_i_shift_amt_2), .A2(ex_block_i_alu_i_shift_amt_3), .ZN(n21894) );
NAND2_X1 U16583 ( .A1(n20830), .A2(n20827), .ZN(n8101) );
NOR2_X1 U16584 ( .A1(n22014), .A2(n15831), .ZN(n21677) );
NOR2_X1 U16585 ( .A1(n22014), .A2(n15836), .ZN(n21671) );
NOR2_X1 U16586 ( .A1(n22014), .A2(n15835), .ZN(n21685) );
NOR2_X1 U16587 ( .A1(n22014), .A2(n15837), .ZN(n21691) );
NOR2_X1 U16588 ( .A1(n16359), .A2(n15838), .ZN(n21780) );
NOR2_X1 U16589 ( .A1(n16359), .A2(n15839), .ZN(n21802) );
NOR2_X1 U16590 ( .A1(n16359), .A2(n15840), .ZN(n21796) );
NOR2_X1 U16591 ( .A1(n16359), .A2(n15841), .ZN(n21738) );
NOR2_X1 U16592 ( .A1(n16359), .A2(n15830), .ZN(n21760) );
NOR2_X1 U16593 ( .A1(n16359), .A2(n15842), .ZN(n21754) );
NOR2_X1 U16594 ( .A1(n16359), .A2(n15834), .ZN(n21842) );
NOR2_X1 U16595 ( .A1(n16359), .A2(n15829), .ZN(n21836) );
NOR2_X1 U16596 ( .A1(n16359), .A2(n15833), .ZN(n21848) );
NOR2_X1 U16597 ( .A1(n22014), .A2(n15854), .ZN(n21710) );
NOR2_X1 U16598 ( .A1(n22014), .A2(n15849), .ZN(n21703) );
NOR2_X1 U16599 ( .A1(n22014), .A2(n15843), .ZN(n21665) );
NOR2_X1 U16600 ( .A1(n16359), .A2(n15850), .ZN(n21770) );
NOR2_X1 U16601 ( .A1(n22014), .A2(n15851), .ZN(n21790) );
NOR2_X1 U16602 ( .A1(n22014), .A2(n15832), .ZN(n21727) );
NOR2_X1 U16603 ( .A1(n22014), .A2(n15852), .ZN(n21748) );
NOR2_X1 U16604 ( .A1(n16359), .A2(n15848), .ZN(n21913) );
NOR2_X1 U16605 ( .A1(n22014), .A2(n15847), .ZN(n21821) );
NOR2_X1 U16606 ( .A1(n22014), .A2(n15855), .ZN(n22003) );
NOR2_X1 U16607 ( .A1(n22014), .A2(n15856), .ZN(n21977) );
NOR2_X1 U16608 ( .A1(n16359), .A2(n15853), .ZN(n21904) );
NOR2_X1 U16609 ( .A1(n16360), .A2(n15832), .ZN(n21912) );
NAND2_X1 U16610 ( .A1(ex_block_i_alu_i_N294), .A2(ex_block_i_alu_i_shift_amt_3), .ZN(n21929) );
NOR2_X1 U16611 ( .A1(n32), .A2(n1416), .ZN(n78) );
NAND2_X1 U16612 ( .A1(n20845), .A2(n20853), .ZN(n9925) );
AND2_X1 U16613 ( .A1(n21929), .A2(n21809), .ZN(n21865) );
NAND2_X1 U16614 ( .A1(ex_block_i_alu_i_N294), .A2(ex_block_i_alu_i_shift_amt_2), .ZN(n21809) );
NAND2_X1 U16615 ( .A1(n7571), .A2(n9918), .ZN(n10044) );
NOR2_X1 U16616 ( .A1(n20939), .A2(n20761), .ZN(n5894) );
NOR2_X1 U16617 ( .A1(n16358), .A2(n15851), .ZN(n21675) );
NOR2_X1 U16618 ( .A1(n16358), .A2(n15838), .ZN(n21683) );
NOR2_X1 U16619 ( .A1(n16358), .A2(n15840), .ZN(n21689) );
NOR2_X1 U16620 ( .A1(n16358), .A2(n15855), .ZN(n21708) );
NOR2_X1 U16621 ( .A1(n16358), .A2(n15850), .ZN(n21701) );
NOR2_X1 U16622 ( .A1(n16351), .A2(n15855), .ZN(n21910) );
NAND2_X1 U16623 ( .A1(n9944), .A2(n20868), .ZN(n7311) );
NOR2_X1 U16624 ( .A1(n22011), .A2(n15839), .ZN(n21669) );
NOR2_X1 U16625 ( .A1(n22011), .A2(n15841), .ZN(n21778) );
NOR2_X1 U16626 ( .A1(n22011), .A2(n15842), .ZN(n21794) );
NOR2_X1 U16627 ( .A1(n22011), .A2(n15834), .ZN(n21736) );
NOR2_X1 U16628 ( .A1(n22011), .A2(n15833), .ZN(n21752) );
NOR2_X1 U16629 ( .A1(n16358), .A2(n15837), .ZN(n21840) );
NOR2_X1 U16630 ( .A1(n16358), .A2(n15835), .ZN(n21825) );
NOR2_X1 U16631 ( .A1(n16358), .A2(n15831), .ZN(n21834) );
NOR2_X1 U16632 ( .A1(n16358), .A2(n15836), .ZN(n21846) );
NOR2_X1 U16633 ( .A1(n16358), .A2(n15844), .ZN(n21663) );
NOR2_X1 U16634 ( .A1(n22011), .A2(n15832), .ZN(n21768) );
NOR2_X1 U16635 ( .A1(n22011), .A2(n15852), .ZN(n21788) );
NOR2_X1 U16636 ( .A1(n22011), .A2(n15848), .ZN(n21725) );
NOR2_X1 U16637 ( .A1(n22011), .A2(n15847), .ZN(n21746) );
NOR2_X1 U16638 ( .A1(n22011), .A2(n15849), .ZN(n21819) );
NOR2_X1 U16639 ( .A1(n22011), .A2(n15856), .ZN(n22001) );
NOR2_X1 U16640 ( .A1(n22011), .A2(n15853), .ZN(n21975) );
NOR2_X1 U16641 ( .A1(n22011), .A2(n15843), .ZN(n21902) );
NOR2_X1 U16642 ( .A1(n15830), .A2(n16358), .ZN(n21800) );
NOR2_X1 U16643 ( .A1(n15829), .A2(n16358), .ZN(n21758) );
NAND2_X1 U16644 ( .A1(n9867), .A2(n9868), .ZN(n9362) );
AND2_X1 U16645 ( .A1(n7571), .A2(n20825), .ZN(n9867) );
NOR2_X1 U16646 ( .A1(n15830), .A2(n16351), .ZN(n21668) );
NOR2_X1 U16647 ( .A1(n15829), .A2(n16351), .ZN(n21799) );
NOR2_X1 U16648 ( .A1(n15831), .A2(n16351), .ZN(n21757) );
NOR2_X1 U16649 ( .A1(n20866), .A2(n15852), .ZN(n21674) );
NOR2_X1 U16650 ( .A1(n20866), .A2(n15841), .ZN(n21682) );
NOR2_X1 U16651 ( .A1(n20866), .A2(n15842), .ZN(n21688) );
NOR2_X1 U16652 ( .A1(n16351), .A2(n15834), .ZN(n21777) );
NOR2_X1 U16653 ( .A1(n16351), .A2(n15833), .ZN(n21793) );
NOR2_X1 U16654 ( .A1(n20866), .A2(n15837), .ZN(n21735) );
NOR2_X1 U16655 ( .A1(n20866), .A2(n15835), .ZN(n21730) );
NOR2_X1 U16656 ( .A1(n20866), .A2(n15836), .ZN(n21751) );
NOR2_X1 U16657 ( .A1(n16351), .A2(n15840), .ZN(n21839) );
NOR2_X1 U16658 ( .A1(n16351), .A2(n15838), .ZN(n21824) );
NOR2_X1 U16659 ( .A1(n16351), .A2(n15851), .ZN(n21833) );
NOR2_X1 U16660 ( .A1(n16351), .A2(n15839), .ZN(n21845) );
NOR2_X1 U16661 ( .A1(n20866), .A2(n15856), .ZN(n21707) );
NOR2_X1 U16662 ( .A1(n20866), .A2(n15832), .ZN(n21700) );
NOR2_X1 U16663 ( .A1(n20866), .A2(n15845), .ZN(n21662) );
NOR2_X1 U16664 ( .A1(n20866), .A2(n15848), .ZN(n21767) );
NOR2_X1 U16665 ( .A1(n20866), .A2(n15847), .ZN(n21787) );
NOR2_X1 U16666 ( .A1(n20866), .A2(n15854), .ZN(n21724) );
NOR2_X1 U16667 ( .A1(n20866), .A2(n15849), .ZN(n21745) );
NOR2_X1 U16668 ( .A1(n20866), .A2(n15850), .ZN(n21818) );
NOR2_X1 U16669 ( .A1(n20866), .A2(n15853), .ZN(n22000) );
NOR2_X1 U16670 ( .A1(n20866), .A2(n15843), .ZN(n21974) );
NOR2_X1 U16671 ( .A1(n20866), .A2(n15844), .ZN(n21901) );
NAND2_X1 U16672 ( .A1(n21673), .A2(n21672), .ZN(n22068) );
NOR2_X1 U16673 ( .A1(n21671), .A2(n21670), .ZN(n21672) );
NOR2_X1 U16674 ( .A1(n21669), .A2(n21668), .ZN(n21673) );
NOR2_X1 U16675 ( .A1(n22015), .A2(n15833), .ZN(n21670) );
NAND2_X1 U16676 ( .A1(n21693), .A2(n21692), .ZN(n21956) );
NOR2_X1 U16677 ( .A1(n21691), .A2(n21690), .ZN(n21692) );
NOR2_X1 U16678 ( .A1(n21689), .A2(n21688), .ZN(n21693) );
NOR2_X1 U16679 ( .A1(n22015), .A2(n15834), .ZN(n21690) );
NAND2_X1 U16680 ( .A1(n21782), .A2(n21781), .ZN(n21895) );
NOR2_X1 U16681 ( .A1(n21780), .A2(n21779), .ZN(n21781) );
NOR2_X1 U16682 ( .A1(n21778), .A2(n21777), .ZN(n21782) );
NOR2_X1 U16683 ( .A1(n16360), .A2(n15835), .ZN(n21779) );
NAND2_X1 U16684 ( .A1(n21804), .A2(n21803), .ZN(n22059) );
NOR2_X1 U16685 ( .A1(n21802), .A2(n21801), .ZN(n21803) );
NOR2_X1 U16686 ( .A1(n21800), .A2(n21799), .ZN(n21804) );
NOR2_X1 U16687 ( .A1(n22015), .A2(n15836), .ZN(n21801) );
NAND2_X1 U16688 ( .A1(n21798), .A2(n21797), .ZN(n21891) );
NOR2_X1 U16689 ( .A1(n21796), .A2(n21795), .ZN(n21797) );
NOR2_X1 U16690 ( .A1(n21794), .A2(n21793), .ZN(n21798) );
NOR2_X1 U16691 ( .A1(n22015), .A2(n15837), .ZN(n21795) );
NAND2_X1 U16692 ( .A1(n21740), .A2(n21739), .ZN(n21885) );
NOR2_X1 U16693 ( .A1(n21738), .A2(n21737), .ZN(n21739) );
NOR2_X1 U16694 ( .A1(n21736), .A2(n21735), .ZN(n21740) );
NOR2_X1 U16695 ( .A1(n16360), .A2(n15838), .ZN(n21737) );
NAND2_X1 U16696 ( .A1(n21762), .A2(n21761), .ZN(n22049) );
NOR2_X1 U16697 ( .A1(n21760), .A2(n21759), .ZN(n21761) );
NOR2_X1 U16698 ( .A1(n21758), .A2(n21757), .ZN(n21762) );
NOR2_X1 U16699 ( .A1(n22015), .A2(n15839), .ZN(n21759) );
NAND2_X1 U16700 ( .A1(n21756), .A2(n21755), .ZN(n21882) );
NOR2_X1 U16701 ( .A1(n21754), .A2(n21753), .ZN(n21755) );
NOR2_X1 U16702 ( .A1(n21752), .A2(n21751), .ZN(n21756) );
NOR2_X1 U16703 ( .A1(n22015), .A2(n15840), .ZN(n21753) );
NAND2_X1 U16704 ( .A1(n21844), .A2(n21843), .ZN(n21962) );
NOR2_X1 U16705 ( .A1(n21842), .A2(n21841), .ZN(n21843) );
NOR2_X1 U16706 ( .A1(n21840), .A2(n21839), .ZN(n21844) );
NOR2_X1 U16707 ( .A1(n16360), .A2(n15841), .ZN(n21841) );
NAND2_X1 U16708 ( .A1(n21838), .A2(n21837), .ZN(n22080) );
NOR2_X1 U16709 ( .A1(n21836), .A2(n21835), .ZN(n21837) );
NOR2_X1 U16710 ( .A1(n21834), .A2(n21833), .ZN(n21838) );
NOR2_X1 U16711 ( .A1(n16360), .A2(n15830), .ZN(n21835) );
NAND2_X1 U16712 ( .A1(n21850), .A2(n21849), .ZN(n22079) );
NOR2_X1 U16713 ( .A1(n21848), .A2(n21847), .ZN(n21849) );
NOR2_X1 U16714 ( .A1(n21846), .A2(n21845), .ZN(n21850) );
NOR2_X1 U16715 ( .A1(n16360), .A2(n15842), .ZN(n21847) );
NAND2_X1 U16716 ( .A1(n21679), .A2(n21678), .ZN(n22069) );
NOR2_X1 U16717 ( .A1(n21677), .A2(n21676), .ZN(n21678) );
NOR2_X1 U16718 ( .A1(n21675), .A2(n21674), .ZN(n21679) );
NOR2_X1 U16719 ( .A1(n15829), .A2(n22015), .ZN(n21676) );
INV_X1 U16720 ( .A(ex_block_i_alu_i_shift_amt_2), .ZN(n20863) );
NOR2_X1 U16721 ( .A1(n20731), .A2(n1708), .ZN(n1730) );
NAND2_X1 U16722 ( .A1(n9944), .A2(n7571), .ZN(n6697) );
INV_X1 U16723 ( .A(n9924), .ZN(n20825) );
NOR2_X1 U16724 ( .A1(n20135), .A2(n10116), .ZN(n10122) );
NOR2_X1 U16725 ( .A1(n21716), .A2(n21715), .ZN(n21717) );
NOR2_X1 U16726 ( .A1(n16360), .A2(n15846), .ZN(n21715) );
NOR2_X1 U16727 ( .A1(n22014), .A2(n16253), .ZN(n21716) );
NOR2_X1 U16728 ( .A1(n22017), .A2(n22016), .ZN(n22018) );
NOR2_X1 U16729 ( .A1(n22015), .A2(n15843), .ZN(n22016) );
NOR2_X1 U16730 ( .A1(n22014), .A2(n15844), .ZN(n22017) );
NOR2_X1 U16731 ( .A1(n21987), .A2(n21986), .ZN(n21988) );
NOR2_X1 U16732 ( .A1(n22015), .A2(n15844), .ZN(n21986) );
NOR2_X1 U16733 ( .A1(n22014), .A2(n15845), .ZN(n21987) );
NOR2_X1 U16734 ( .A1(n21919), .A2(n21918), .ZN(n21920) );
NOR2_X1 U16735 ( .A1(n22015), .A2(n15845), .ZN(n21918) );
NOR2_X1 U16736 ( .A1(n22014), .A2(n15846), .ZN(n21919) );
NAND2_X1 U16737 ( .A1(n21915), .A2(n21914), .ZN(n22039) );
NOR2_X1 U16738 ( .A1(n21911), .A2(n21910), .ZN(n21915) );
NOR2_X1 U16739 ( .A1(n21913), .A2(n21912), .ZN(n21914) );
NOR2_X1 U16740 ( .A1(n22011), .A2(n15854), .ZN(n21911) );
NOR2_X1 U16741 ( .A1(n10032), .A2(n10033), .ZN(n10031) );
NAND2_X1 U16742 ( .A1(n10036), .A2(n20861), .ZN(n10032) );
NAND2_X1 U16743 ( .A1(n10034), .A2(n10035), .ZN(n10033) );
NAND2_X1 U16744 ( .A1(n20827), .A2(n20838), .ZN(n10036) );
NOR2_X1 U16745 ( .A1(n1383), .A2(n1384), .ZN(n1382) );
NAND2_X1 U16746 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
NOR2_X1 U16747 ( .A1(n1335), .A2(n16247), .ZN(n1383) );
NAND2_X1 U16748 ( .A1(n1387), .A2(n20759), .ZN(n1386) );
NAND2_X1 U16749 ( .A1(n9938), .A2(n7571), .ZN(n8584) );
NOR2_X1 U16750 ( .A1(n1565), .A2(n15797), .ZN(n6513) );
INV_X1 U16751 ( .A(ex_block_i_alu_i_shift_operand_31), .ZN(n20134) );
NOR2_X1 U16752 ( .A1(n21714), .A2(n21713), .ZN(n21718) );
AND2_X1 U16753 ( .A1(ex_block_i_alu_i_shift_operand_0), .A2(n21773), .ZN(n21713) );
NOR2_X1 U16754 ( .A1(n22011), .A2(n16256), .ZN(n21714) );
NAND2_X1 U16755 ( .A1(n5797), .A2(n5798), .ZN(ex_block_i_alu_i_shift_operand_0) );
NOR2_X1 U16756 ( .A1(n22013), .A2(n22012), .ZN(n22019) );
NOR2_X1 U16757 ( .A1(n22011), .A2(n15845), .ZN(n22013) );
NOR2_X1 U16758 ( .A1(n20866), .A2(n15846), .ZN(n22012) );
NOR2_X1 U16759 ( .A1(n21985), .A2(n21984), .ZN(n21989) );
NOR2_X1 U16760 ( .A1(n22011), .A2(n15846), .ZN(n21985) );
NOR2_X1 U16761 ( .A1(n16351), .A2(n16253), .ZN(n21984) );
NOR2_X1 U16762 ( .A1(n21917), .A2(n21916), .ZN(n21921) );
NOR2_X1 U16763 ( .A1(n22011), .A2(n16253), .ZN(n21917) );
NOR2_X1 U16764 ( .A1(n16351), .A2(n16256), .ZN(n21916) );
NAND2_X1 U16765 ( .A1(n20859), .A2(n20853), .ZN(n9844) );
INV_X1 U16766 ( .A(ex_block_i_alu_i_shift_amt_3), .ZN(n20856) );
INV_X1 U16767 ( .A(n7657), .ZN(n20885) );
NAND2_X1 U16768 ( .A1(n10019), .A2(n1432), .ZN(n8122) );
NOR2_X1 U16769 ( .A1(n20833), .A2(n20835), .ZN(n10019) );
NAND2_X1 U16770 ( .A1(n78), .A2(n260), .ZN(n259) );
NAND2_X1 U16771 ( .A1(n7638), .A2(n7639), .ZN(n4049) );
NAND2_X1 U16772 ( .A1(n20985), .A2(n7659), .ZN(n7638) );
NAND2_X1 U16773 ( .A1(n7581), .A2(n7640), .ZN(n7639) );
NAND2_X1 U16774 ( .A1(n7660), .A2(n7661), .ZN(n7659) );
NAND2_X1 U16775 ( .A1(n21775), .A2(n21774), .ZN(n21863) );
NAND2_X1 U16776 ( .A1(ex_block_i_alu_i_shift_operand_31), .A2(n21773), .ZN(n21775) );
NAND2_X1 U16777 ( .A1(ex_block_i_alu_i_N294), .A2(n16351), .ZN(n21774) );
NAND2_X1 U16778 ( .A1(n21733), .A2(n21732), .ZN(n21855) );
NAND2_X1 U16779 ( .A1(ex_block_i_alu_i_N294), .A2(ex_block_i_alu_i_shift_amt_1), .ZN(n21732) );
NOR2_X1 U16780 ( .A1(n21731), .A2(n21730), .ZN(n21733) );
NOR2_X1 U16781 ( .A1(n22011), .A2(n20134), .ZN(n21731) );
NAND2_X1 U16782 ( .A1(n21705), .A2(n21704), .ZN(n22030) );
NOR2_X1 U16783 ( .A1(n21703), .A2(n21702), .ZN(n21704) );
NOR2_X1 U16784 ( .A1(n21701), .A2(n21700), .ZN(n21705) );
NOR2_X1 U16785 ( .A1(n16360), .A2(n15847), .ZN(n21702) );
NAND2_X1 U16786 ( .A1(n21712), .A2(n21711), .ZN(n22029) );
NOR2_X1 U16787 ( .A1(n21710), .A2(n21709), .ZN(n21711) );
NOR2_X1 U16788 ( .A1(n21708), .A2(n21707), .ZN(n21712) );
NOR2_X1 U16789 ( .A1(n16360), .A2(n15848), .ZN(n21709) );
NAND2_X1 U16790 ( .A1(n21772), .A2(n21771), .ZN(n22010) );
NOR2_X1 U16791 ( .A1(n21770), .A2(n21769), .ZN(n21771) );
NOR2_X1 U16792 ( .A1(n21768), .A2(n21767), .ZN(n21772) );
NOR2_X1 U16793 ( .A1(n22015), .A2(n15849), .ZN(n21769) );
NAND2_X1 U16794 ( .A1(n21792), .A2(n21791), .ZN(n22060) );
NOR2_X1 U16795 ( .A1(n21790), .A2(n21789), .ZN(n21791) );
NOR2_X1 U16796 ( .A1(n21788), .A2(n21787), .ZN(n21792) );
NOR2_X1 U16797 ( .A1(n22015), .A2(n15831), .ZN(n21789) );
NAND2_X1 U16798 ( .A1(n21729), .A2(n21728), .ZN(n21983) );
NOR2_X1 U16799 ( .A1(n21727), .A2(n21726), .ZN(n21728) );
NOR2_X1 U16800 ( .A1(n21725), .A2(n21724), .ZN(n21729) );
NOR2_X1 U16801 ( .A1(n16360), .A2(n15850), .ZN(n21726) );
NAND2_X1 U16802 ( .A1(n21750), .A2(n21749), .ZN(n22050) );
NOR2_X1 U16803 ( .A1(n21748), .A2(n21747), .ZN(n21749) );
NOR2_X1 U16804 ( .A1(n21746), .A2(n21745), .ZN(n21750) );
NOR2_X1 U16805 ( .A1(n16360), .A2(n15851), .ZN(n21747) );
NAND2_X1 U16806 ( .A1(n21823), .A2(n21822), .ZN(n22040) );
NOR2_X1 U16807 ( .A1(n21821), .A2(n21820), .ZN(n21822) );
NOR2_X1 U16808 ( .A1(n21819), .A2(n21818), .ZN(n21823) );
NOR2_X1 U16809 ( .A1(n22015), .A2(n15852), .ZN(n21820) );
AND2_X1 U16810 ( .A1(n21667), .A2(n21666), .ZN(n22025) );
NOR2_X1 U16811 ( .A1(n21665), .A2(n21664), .ZN(n21666) );
NOR2_X1 U16812 ( .A1(n21663), .A2(n21662), .ZN(n21667) );
NOR2_X1 U16813 ( .A1(n16360), .A2(n15853), .ZN(n21664) );
AND2_X1 U16814 ( .A1(n22005), .A2(n22004), .ZN(n22055) );
NOR2_X1 U16815 ( .A1(n22003), .A2(n22002), .ZN(n22004) );
NOR2_X1 U16816 ( .A1(n22001), .A2(n22000), .ZN(n22005) );
NOR2_X1 U16817 ( .A1(n22015), .A2(n15854), .ZN(n22002) );
AND2_X1 U16818 ( .A1(n21979), .A2(n21978), .ZN(n22045) );
NOR2_X1 U16819 ( .A1(n21977), .A2(n21976), .ZN(n21978) );
NOR2_X1 U16820 ( .A1(n21975), .A2(n21974), .ZN(n21979) );
NOR2_X1 U16821 ( .A1(n22015), .A2(n15855), .ZN(n21976) );
AND2_X1 U16822 ( .A1(n21906), .A2(n21905), .ZN(n22035) );
NOR2_X1 U16823 ( .A1(n21904), .A2(n21903), .ZN(n21905) );
NOR2_X1 U16824 ( .A1(n21902), .A2(n21901), .ZN(n21906) );
NOR2_X1 U16825 ( .A1(n16360), .A2(n15856), .ZN(n21903) );
AND2_X1 U16826 ( .A1(n21229), .A2(n21228), .ZN(n21230) );
NOR2_X1 U16827 ( .A1(n21229), .A2(n21228), .ZN(n21231) );
NAND2_X1 U16828 ( .A1(n21227), .A2(n21226), .ZN(n21228) );
INV_X1 U16829 ( .A(n10115), .ZN(n20135) );
NAND2_X1 U16830 ( .A1(n9970), .A2(n20864), .ZN(n10045) );
NAND2_X1 U16831 ( .A1(n9906), .A2(n9907), .ZN(n8567) );
NOR2_X1 U16832 ( .A1(n9908), .A2(n8312), .ZN(n9906) );
NAND2_X1 U16833 ( .A1(n9914), .A2(n9907), .ZN(n8572) );
NOR2_X1 U16834 ( .A1(n9841), .A2(n8312), .ZN(n9914) );
NAND2_X1 U16835 ( .A1(n32), .A2(n16335), .ZN(rf_we_wb_o) );
NAND2_X1 U16836 ( .A1(ex_block_i_alu_i_shift_amt_0), .A2(n20867), .ZN(n22011) );
INV_X1 U16837 ( .A(n7678), .ZN(n20886) );
INV_X1 U16838 ( .A(ex_block_i_alu_i_shift_amt_1), .ZN(n20867) );
NAND2_X1 U16839 ( .A1(n20832), .A2(n5245), .ZN(n10018) );
AND2_X1 U16840 ( .A1(n21872), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n21698) );
AND2_X1 U16841 ( .A1(n21997), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n21866) );
AND2_X1 U16842 ( .A1(n21995), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n21857) );
AND2_X1 U16843 ( .A1(n21972), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n21831) );
AND2_X1 U16844 ( .A1(n21970), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n21812) );
AND2_X1 U16845 ( .A1(n21968), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n21785) );
AND2_X1 U16846 ( .A1(n21966), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n21743) );
AND2_X1 U16847 ( .A1(n22075), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n22076) );
AND2_X1 U16848 ( .A1(n22065), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n22066) );
AND2_X1 U16849 ( .A1(n22056), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n22057) );
AND2_X1 U16850 ( .A1(n22046), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n22047) );
AND2_X1 U16851 ( .A1(n22036), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n22037) );
AND2_X1 U16852 ( .A1(n22026), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n22027) );
AND2_X1 U16853 ( .A1(n22006), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n22007) );
AND2_X1 U16854 ( .A1(n21980), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n21981) );
AND2_X1 U16855 ( .A1(n21907), .A2(ex_block_i_alu_i_shift_amt_4), .ZN(n21908) );
INV_X1 U16856 ( .A(n7684), .ZN(n20890) );
INV_X1 U16857 ( .A(ex_block_i_alu_i_adder_in_a_3), .ZN(n20750) );
INV_X1 U16858 ( .A(ex_block_i_alu_i_adder_in_a_4), .ZN(n20744) );
INV_X1 U16859 ( .A(ex_block_i_alu_i_adder_in_a_5), .ZN(n20739) );
INV_X1 U16860 ( .A(ex_block_i_alu_i_adder_in_a_6), .ZN(n20733) );
INV_X1 U16861 ( .A(ex_block_i_alu_i_adder_in_a_7), .ZN(n20728) );
INV_X1 U16862 ( .A(ex_block_i_alu_i_adder_in_a_8), .ZN(n20722) );
INV_X1 U16863 ( .A(ex_block_i_alu_i_adder_in_a_9), .ZN(n20717) );
INV_X1 U16864 ( .A(ex_block_i_alu_i_adder_in_a_10), .ZN(n20713) );
INV_X1 U16865 ( .A(ex_block_i_alu_i_adder_in_a_2), .ZN(n20754) );
INV_X1 U16866 ( .A(ex_block_i_alu_i_adder_in_a_11), .ZN(n20709) );
INV_X1 U16867 ( .A(ex_block_i_alu_i_adder_in_a_12), .ZN(n20705) );
INV_X1 U16868 ( .A(ex_block_i_alu_i_adder_in_a_13), .ZN(n20701) );
INV_X1 U16869 ( .A(ex_block_i_alu_i_adder_in_a_14), .ZN(n20697) );
INV_X1 U16870 ( .A(ex_block_i_alu_i_adder_in_a_15), .ZN(n20693) );
INV_X1 U16871 ( .A(ex_block_i_alu_i_adder_in_a_16), .ZN(n20689) );
INV_X1 U16872 ( .A(ex_block_i_alu_i_adder_in_a_17), .ZN(n20685) );
INV_X1 U16873 ( .A(ex_block_i_alu_i_adder_in_a_18), .ZN(n20678) );
INV_X1 U16874 ( .A(ex_block_i_alu_i_adder_in_a_19), .ZN(n20644) );
INV_X1 U16875 ( .A(ex_block_i_alu_i_adder_in_a_20), .ZN(n20606) );
INV_X1 U16876 ( .A(ex_block_i_alu_i_adder_in_a_21), .ZN(n20566) );
INV_X1 U16877 ( .A(ex_block_i_alu_i_adder_in_a_22), .ZN(n20526) );
INV_X1 U16878 ( .A(ex_block_i_alu_i_adder_in_a_23), .ZN(n20486) );
INV_X1 U16879 ( .A(ex_block_i_alu_i_adder_in_a_24), .ZN(n20446) );
INV_X1 U16880 ( .A(ex_block_i_alu_i_adder_in_a_25), .ZN(n20406) );
INV_X1 U16881 ( .A(ex_block_i_alu_i_adder_in_a_26), .ZN(n20367) );
INV_X1 U16882 ( .A(ex_block_i_alu_i_adder_in_a_27), .ZN(n20328) );
INV_X1 U16883 ( .A(ex_block_i_alu_i_adder_in_a_28), .ZN(n20289) );
INV_X1 U16884 ( .A(ex_block_i_alu_i_adder_in_a_29), .ZN(n20250) );
INV_X1 U16885 ( .A(ex_block_i_alu_i_adder_in_a_30), .ZN(n20212) );
INV_X1 U16886 ( .A(ex_block_i_alu_i_adder_in_a_31), .ZN(n20174) );
NAND2_X1 U16887 ( .A1(ex_block_i_alu_i_adder_in_b_20), .A2(n20606), .ZN(n21140) );
NAND2_X1 U16888 ( .A1(ex_block_i_alu_i_adder_in_b_21), .A2(n20566), .ZN(n21149) );
NAND2_X1 U16889 ( .A1(ex_block_i_alu_i_adder_in_b_22), .A2(n20526), .ZN(n21158) );
NAND2_X1 U16890 ( .A1(ex_block_i_alu_i_adder_in_b_23), .A2(n20486), .ZN(n21167) );
NAND2_X1 U16891 ( .A1(ex_block_i_alu_i_adder_in_b_24), .A2(n20446), .ZN(n21176) );
NAND2_X1 U16892 ( .A1(ex_block_i_alu_i_adder_in_b_25), .A2(n20406), .ZN(n21185) );
NAND2_X1 U16893 ( .A1(ex_block_i_alu_i_adder_in_b_26), .A2(n20367), .ZN(n21194) );
NAND2_X1 U16894 ( .A1(ex_block_i_alu_i_adder_in_b_27), .A2(n20328), .ZN(n21203) );
NAND2_X1 U16895 ( .A1(ex_block_i_alu_i_adder_in_b_28), .A2(n20289), .ZN(n21212) );
NAND2_X1 U16896 ( .A1(ex_block_i_alu_i_adder_in_b_29), .A2(n20250), .ZN(n21221) );
NAND2_X1 U16897 ( .A1(ex_block_i_alu_i_adder_in_b_30), .A2(n20212), .ZN(n21236) );
NAND2_X1 U16898 ( .A1(ex_block_i_alu_i_adder_in_b_31), .A2(n20174), .ZN(n21245) );
NAND2_X1 U16899 ( .A1(ex_block_i_alu_i_adder_in_b_13), .A2(n20701), .ZN(n21072) );
NAND2_X1 U16900 ( .A1(ex_block_i_alu_i_adder_in_b_14), .A2(n20697), .ZN(n21081) );
NAND2_X1 U16901 ( .A1(ex_block_i_alu_i_adder_in_b_15), .A2(n20693), .ZN(n21090) );
NAND2_X1 U16902 ( .A1(ex_block_i_alu_i_adder_in_b_16), .A2(n20689), .ZN(n21099) );
NAND2_X1 U16903 ( .A1(ex_block_i_alu_i_adder_in_b_17), .A2(n20685), .ZN(n21108) );
NAND2_X1 U16904 ( .A1(ex_block_i_alu_i_adder_in_b_18), .A2(n20678), .ZN(n21117) );
NAND2_X1 U16905 ( .A1(ex_block_i_alu_i_adder_in_b_19), .A2(n20644), .ZN(n21126) );
OR2_X1 U16906 ( .A1(n20893), .A2(n7619), .ZN(n7618) );
NAND2_X1 U16907 ( .A1(n20940), .A2(n20944), .ZN(n6304) );
NAND2_X1 U16908 ( .A1(n6305), .A2(n20945), .ZN(n6303) );
AND2_X1 U16909 ( .A1(n6306), .A2(ex_block_i_alu_i_shift_operand_31), .ZN(n6305) );
OR2_X1 U16910 ( .A1(n20697), .A2(ex_block_i_alu_i_adder_in_b_14), .ZN(n21082) );
OR2_X1 U16911 ( .A1(n20685), .A2(ex_block_i_alu_i_adder_in_b_17), .ZN(n21109) );
OR2_X1 U16912 ( .A1(n20678), .A2(ex_block_i_alu_i_adder_in_b_18), .ZN(n21118) );
OR2_X1 U16913 ( .A1(n20566), .A2(ex_block_i_alu_i_adder_in_b_21), .ZN(n21150) );
OR2_X1 U16914 ( .A1(n20446), .A2(ex_block_i_alu_i_adder_in_b_24), .ZN(n21177) );
OR2_X1 U16915 ( .A1(n20328), .A2(ex_block_i_alu_i_adder_in_b_27), .ZN(n21204) );
OR2_X1 U16916 ( .A1(n20289), .A2(ex_block_i_alu_i_adder_in_b_28), .ZN(n21213) );
OR2_X1 U16917 ( .A1(n20174), .A2(ex_block_i_alu_i_adder_in_b_31), .ZN(n21246) );
OR2_X1 U16918 ( .A1(n20701), .A2(ex_block_i_alu_i_adder_in_b_13), .ZN(n21073) );
OR2_X1 U16919 ( .A1(n20693), .A2(ex_block_i_alu_i_adder_in_b_15), .ZN(n21091) );
OR2_X1 U16920 ( .A1(n20689), .A2(ex_block_i_alu_i_adder_in_b_16), .ZN(n21100) );
OR2_X1 U16921 ( .A1(n20644), .A2(ex_block_i_alu_i_adder_in_b_19), .ZN(n21127) );
OR2_X1 U16922 ( .A1(n20606), .A2(ex_block_i_alu_i_adder_in_b_20), .ZN(n21141) );
OR2_X1 U16923 ( .A1(n20526), .A2(ex_block_i_alu_i_adder_in_b_22), .ZN(n21159) );
OR2_X1 U16924 ( .A1(n20486), .A2(ex_block_i_alu_i_adder_in_b_23), .ZN(n21168) );
OR2_X1 U16925 ( .A1(n20406), .A2(ex_block_i_alu_i_adder_in_b_25), .ZN(n21186) );
OR2_X1 U16926 ( .A1(n20367), .A2(ex_block_i_alu_i_adder_in_b_26), .ZN(n21195) );
OR2_X1 U16927 ( .A1(n20250), .A2(ex_block_i_alu_i_adder_in_b_29), .ZN(n21222) );
OR2_X1 U16928 ( .A1(n20212), .A2(ex_block_i_alu_i_adder_in_b_30), .ZN(n21237) );
NAND2_X1 U16929 ( .A1(n21135), .A2(n21134), .ZN(alu_adder_result_ex_0) );
NAND2_X1 U16930 ( .A1(n21133), .A2(n20758), .ZN(n21135) );
OR2_X1 U16931 ( .A1(n21133), .A2(n20758), .ZN(n21134) );
NAND2_X1 U16932 ( .A1(n21132), .A2(n21131), .ZN(n21133) );
NAND2_X1 U16933 ( .A1(ex_block_i_alu_i_shift_amt_0), .A2(ex_block_i_alu_i_shift_amt_1), .ZN(n22015) );
OR2_X1 U16934 ( .A1(n20867), .A2(ex_block_i_alu_i_shift_amt_0), .ZN(n22014) );
NAND2_X1 U16935 ( .A1(n1065), .A2(n1039), .ZN(n378) );
NOR2_X1 U16936 ( .A1(n1058), .A2(n16335), .ZN(n1065) );
NAND2_X1 U16937 ( .A1(n1364), .A2(n19967), .ZN(n45) );
NOR2_X1 U16938 ( .A1(n1373), .A2(n1058), .ZN(n1364) );
NOR2_X1 U16939 ( .A1(n21017), .A2(n1039), .ZN(n1373) );
BUF_X1 U16940 ( .A(n44), .Z(n16477) );
INV_X1 U16941 ( .A(n33), .ZN(n19967) );
NOR2_X1 U16942 ( .A1(n20871), .A2(n1317), .ZN(n1396) );
NOR2_X1 U16943 ( .A1(n20871), .A2(n1319), .ZN(n1387) );
INV_X1 U16944 ( .A(n363), .ZN(n19966) );
INV_X1 U16945 ( .A(n16399), .ZN(n16400) );
INV_X1 U16946 ( .A(n16399), .ZN(n16401) );
NAND2_X1 U16947 ( .A1(n21001), .A2(n5091), .ZN(n5911) );
NAND2_X1 U16948 ( .A1(n6719), .A2(n7023), .ZN(n6711) );
BUF_X1 U16949 ( .A(n4291), .Z(n16419) );
INV_X1 U16950 ( .A(n6793), .ZN(n20876) );
AND2_X1 U16951 ( .A1(n4417), .A2(n4918), .ZN(n4447) );
BUF_X1 U16952 ( .A(n6708), .Z(n16403) );
INV_X1 U16953 ( .A(n5374), .ZN(n20906) );
INV_X1 U16954 ( .A(n6796), .ZN(n20875) );
OR2_X1 U16955 ( .A1(n5272), .A2(n5736), .ZN(n5674) );
BUF_X1 U16956 ( .A(n6238), .Z(n16408) );
BUF_X1 U16957 ( .A(n4272), .Z(n16424) );
BUF_X1 U16958 ( .A(n4288), .Z(n16420) );
BUF_X1 U16959 ( .A(n7872), .Z(n16389) );
AND2_X1 U16960 ( .A1(n4447), .A2(n4917), .ZN(n4270) );
NAND2_X1 U16961 ( .A1(n1422), .A2(n1423), .ZN(n4917) );
NAND2_X1 U16962 ( .A1(n20956), .A2(n10156), .ZN(n5910) );
INV_X1 U16963 ( .A(n5916), .ZN(n20959) );
INV_X1 U16964 ( .A(n5917), .ZN(n20960) );
NOR2_X1 U16965 ( .A1(n1435), .A2(n1416), .ZN(n1432) );
BUF_X1 U16966 ( .A(n4287), .Z(n16421) );
BUF_X1 U16967 ( .A(n3263), .Z(n16433) );
BUF_X1 U16968 ( .A(n7875), .Z(n16388) );
NAND2_X1 U16969 ( .A1(n20948), .A2(n20949), .ZN(n8773) );
BUF_X1 U16970 ( .A(n5268), .Z(n16418) );
INV_X1 U16971 ( .A(n7084), .ZN(n19983) );
NOR2_X1 U16972 ( .A1(n2058), .A2(n2410), .ZN(n2026) );
BUF_X1 U16973 ( .A(n20917), .Z(n16353) );
NOR2_X1 U16974 ( .A1(n2655), .A2(n2557), .ZN(n2332) );
BUF_X1 U16975 ( .A(n3130), .Z(n16435) );
NOR2_X1 U16976 ( .A1(n2715), .A2(n2058), .ZN(n2055) );
NOR2_X1 U16977 ( .A1(n19941), .A2(n2715), .ZN(n2049) );
NAND2_X1 U16978 ( .A1(n21017), .A2(n21016), .ZN(n72) );
INV_X1 U16979 ( .A(n6306), .ZN(n20952) );
NOR2_X1 U16980 ( .A1(n20984), .A2(n20929), .ZN(n4005) );
NOR2_X1 U16981 ( .A1(n2557), .A2(n2058), .ZN(n2029) );
NOR2_X1 U16982 ( .A1(n16399), .A2(n5147), .ZN(n7019) );
AND2_X1 U16983 ( .A1(n21014), .A2(n1325), .ZN(n70) );
OR2_X1 U16984 ( .A1(n1039), .A2(n21017), .ZN(n1325) );
NAND2_X1 U16985 ( .A1(n2142), .A2(n2302), .ZN(n2222) );
NAND2_X1 U16986 ( .A1(n2303), .A2(n2204), .ZN(n2302) );
NAND2_X1 U16987 ( .A1(n4004), .A2(n4005), .ZN(n3776) );
NOR2_X1 U16988 ( .A1(n20928), .A2(n3777), .ZN(n4004) );
NOR2_X1 U16989 ( .A1(n5826), .A2(n5091), .ZN(n5904) );
NAND2_X1 U16990 ( .A1(n20986), .A2(n5125), .ZN(n7041) );
NAND2_X1 U16991 ( .A1(n8824), .A2(n8825), .ZN(n7037) );
NAND2_X1 U16992 ( .A1(n8826), .A2(n20745), .ZN(n8825) );
NAND2_X1 U16993 ( .A1(n323), .A2(n16418), .ZN(n8824) );
INV_X1 U16994 ( .A(n323), .ZN(n20745) );
NAND2_X1 U16995 ( .A1(n7569), .A2(n7718), .ZN(n7577) );
NAND2_X1 U16996 ( .A1(n7032), .A2(n7719), .ZN(n7718) );
NOR2_X1 U16997 ( .A1(n10273), .A2(data_we_o), .ZN(n6509) );
NOR2_X1 U16998 ( .A1(n1435), .A2(n1596), .ZN(n10273) );
INV_X1 U16999 ( .A(n7069), .ZN(n19789) );
INV_X1 U17000 ( .A(n7203), .ZN(n19807) );
INV_X1 U17001 ( .A(n7068), .ZN(n19787) );
NOR2_X1 U17002 ( .A1(n16454), .A2(n1447), .ZN(n3567) );
INV_X1 U17003 ( .A(n7237), .ZN(n19781) );
INV_X1 U17004 ( .A(n6792), .ZN(n19749) );
INV_X1 U17005 ( .A(n7243), .ZN(n19785) );
INV_X1 U17006 ( .A(n7185), .ZN(n19797) );
INV_X1 U17007 ( .A(n7240), .ZN(n19783) );
INV_X1 U17008 ( .A(n7250), .ZN(n19791) );
INV_X1 U17009 ( .A(n7179), .ZN(n19793) );
INV_X1 U17010 ( .A(n7182), .ZN(n19795) );
NOR2_X1 U17011 ( .A1(n2409), .A2(n2058), .ZN(n2363) );
INV_X1 U17012 ( .A(n7253), .ZN(n19811) );
NOR2_X1 U17013 ( .A1(n20961), .A2(n20962), .ZN(n1423) );
INV_X1 U17014 ( .A(n897), .ZN(n21012) );
INV_X1 U17015 ( .A(n898), .ZN(n21015) );
NOR2_X1 U17016 ( .A1(n2715), .A2(n19940), .ZN(n2397) );
INV_X1 U17017 ( .A(n6896), .ZN(n19769) );
INV_X1 U17018 ( .A(n6943), .ZN(n19777) );
AND2_X1 U17019 ( .A1(n8129), .A2(n8130), .ZN(n8128) );
NOR2_X1 U17020 ( .A1(n20841), .A2(n8115), .ZN(n8130) );
INV_X1 U17021 ( .A(n6842), .ZN(n19757) );
INV_X1 U17022 ( .A(n6851), .ZN(n19759) );
INV_X1 U17023 ( .A(n6860), .ZN(n19761) );
INV_X1 U17024 ( .A(n6869), .ZN(n19763) );
INV_X1 U17025 ( .A(n6878), .ZN(n19765) );
INV_X1 U17026 ( .A(n6887), .ZN(n19767) );
INV_X1 U17027 ( .A(n6905), .ZN(n19771) );
INV_X1 U17028 ( .A(n6925), .ZN(n19773) );
INV_X1 U17029 ( .A(n6934), .ZN(n19775) );
INV_X1 U17030 ( .A(n6952), .ZN(n19779) );
INV_X1 U17031 ( .A(n6833), .ZN(n19755) );
INV_X1 U17032 ( .A(n6803), .ZN(n19751) );
INV_X1 U17033 ( .A(n6824), .ZN(n19753) );
INV_X1 U17034 ( .A(n7191), .ZN(n19801) );
INV_X1 U17035 ( .A(n7188), .ZN(n19799) );
INV_X1 U17036 ( .A(n2270), .ZN(n19940) );
NAND2_X1 U17037 ( .A1(n16451), .A2(n2060), .ZN(n2471) );
NOR2_X1 U17038 ( .A1(n16400), .A2(n7580), .ZN(n7569) );
INV_X1 U17039 ( .A(n4051), .ZN(n20991) );
NOR2_X1 U17040 ( .A1(n2303), .A2(n19881), .ZN(n2339) );
NOR2_X1 U17041 ( .A1(n2204), .A2(n19881), .ZN(n2178) );
NAND2_X1 U17042 ( .A1(n2766), .A2(n19907), .ZN(n2557) );
NOR2_X1 U17043 ( .A1(n19910), .A2(n19912), .ZN(n2766) );
NAND2_X1 U17044 ( .A1(n8778), .A2(n8779), .ZN(n7194) );
NAND2_X1 U17045 ( .A1(n8780), .A2(n20740), .ZN(n8779) );
NAND2_X1 U17046 ( .A1(n282), .A2(n16418), .ZN(n8778) );
INV_X1 U17047 ( .A(n282), .ZN(n20740) );
NAND2_X1 U17048 ( .A1(n9387), .A2(n9388), .ZN(n7226) );
NAND2_X1 U17049 ( .A1(n9389), .A2(n20755), .ZN(n9388) );
NAND2_X1 U17050 ( .A1(n883), .A2(n5268), .ZN(n9387) );
INV_X1 U17051 ( .A(n883), .ZN(n20755) );
NOR2_X1 U17052 ( .A1(n7067), .A2(n7052), .ZN(n7059) );
NOR2_X1 U17053 ( .A1(n7068), .A2(n7069), .ZN(n7067) );
NAND2_X1 U17054 ( .A1(n16400), .A2(n20880), .ZN(n7323) );
NOR2_X1 U17055 ( .A1(n2456), .A2(n19914), .ZN(n2047) );
NOR2_X1 U17056 ( .A1(n10275), .A2(n10266), .ZN(n5108) );
AND2_X1 U17057 ( .A1(n10276), .A2(n10277), .ZN(n10275) );
NAND2_X1 U17058 ( .A1(n20920), .A2(n20912), .ZN(n10277) );
NOR2_X1 U17059 ( .A1(n1395), .A2(n20944), .ZN(n10117) );
NAND2_X1 U17060 ( .A1(n4417), .A2(n20962), .ZN(n4412) );
NOR2_X1 U17061 ( .A1(n22100), .A2(n22089), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_16) );
NOR2_X1 U17062 ( .A1(n22100), .A2(n22092), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_24) );
NOR2_X1 U17063 ( .A1(n20945), .A2(n6231), .ZN(n6309) );
NOR2_X1 U17064 ( .A1(n2538), .A2(n2539), .ZN(n2352) );
AND2_X1 U17065 ( .A1(n2047), .A2(n2048), .ZN(n2538) );
NOR2_X1 U17066 ( .A1(n5129), .A2(n20989), .ZN(n5143) );
NOR2_X1 U17067 ( .A1(n20986), .A2(n20991), .ZN(n5225) );
INV_X1 U17068 ( .A(n1435), .ZN(n20912) );
INV_X1 U17069 ( .A(n2409), .ZN(n19904) );
NOR2_X1 U17070 ( .A1(n19929), .A2(n2470), .ZN(n2686) );
NOR2_X1 U17071 ( .A1(n19917), .A2(n19919), .ZN(n2675) );
NOR2_X1 U17072 ( .A1(n16461), .A2(n1687), .ZN(n1657) );
INV_X1 U17073 ( .A(n5147), .ZN(n20985) );
INV_X1 U17074 ( .A(n2715), .ZN(n19906) );
INV_X1 U17075 ( .A(n4998), .ZN(n21008) );
NAND2_X1 U17076 ( .A1(n5540), .A2(n20919), .ZN(n4411) );
NOR2_X1 U17077 ( .A1(n22100), .A2(n22096), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_0) );
NOR2_X1 U17078 ( .A1(n22100), .A2(n22099), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_8) );
NAND2_X1 U17079 ( .A1(n19912), .A2(n19891), .ZN(n2113) );
NAND2_X1 U17080 ( .A1(n10517), .A2(n10145), .ZN(n10501) );
NOR2_X1 U17081 ( .A1(n10141), .A2(n1687), .ZN(n10517) );
NAND2_X1 U17082 ( .A1(n2172), .A2(n2142), .ZN(n2156) );
NAND2_X1 U17083 ( .A1(n2697), .A2(n2349), .ZN(n2184) );
NOR2_X1 U17084 ( .A1(n3586), .A2(n3587), .ZN(n1885) );
AND2_X1 U17085 ( .A1(n3588), .A2(n3589), .ZN(n3587) );
NOR2_X1 U17086 ( .A1(n16449), .A2(n3592), .ZN(n3588) );
NOR2_X1 U17087 ( .A1(n3590), .A2(n3591), .ZN(n3589) );
NOR2_X1 U17088 ( .A1(n1435), .A2(n20822), .ZN(n5242) );
NAND2_X1 U17089 ( .A1(n2049), .A2(n2456), .ZN(n2182) );
NAND2_X1 U17090 ( .A1(n8096), .A2(n7082), .ZN(n8083) );
NOR2_X1 U17091 ( .A1(n7078), .A2(n7084), .ZN(n8096) );
AND2_X1 U17092 ( .A1(n2619), .A2(n2582), .ZN(n2152) );
NAND2_X1 U17093 ( .A1(n2112), .A2(n19890), .ZN(n2619) );
INV_X1 U17094 ( .A(n1606), .ZN(n16461) );
INV_X1 U17095 ( .A(n8600), .ZN(n16366) );
INV_X1 U17096 ( .A(n2756), .ZN(n20903) );
NOR2_X1 U17097 ( .A1(n1446), .A2(n20747), .ZN(n21384) );
NOR2_X1 U17098 ( .A1(n20997), .A2(n20996), .ZN(n1518) );
NOR2_X1 U17099 ( .A1(n6234), .A2(n20952), .ZN(n1411) );
NAND2_X1 U17100 ( .A1(n2522), .A2(n2410), .ZN(n2453) );
INV_X1 U17101 ( .A(n5011), .ZN(n21009) );
NOR2_X1 U17102 ( .A1(n8118), .A2(n7084), .ZN(n8129) );
NOR2_X1 U17103 ( .A1(n2594), .A2(n19881), .ZN(n2593) );
NOR2_X1 U17104 ( .A1(n2595), .A2(n2596), .ZN(n2594) );
NAND2_X1 U17105 ( .A1(n2600), .A2(n2601), .ZN(n2595) );
NAND2_X1 U17106 ( .A1(n19892), .A2(n2598), .ZN(n2596) );
NOR2_X1 U17107 ( .A1(n16399), .A2(n20880), .ZN(n7319) );
INV_X1 U17108 ( .A(n6231), .ZN(n20944) );
NAND2_X1 U17109 ( .A1(n2113), .A2(n2697), .ZN(n2269) );
INV_X1 U17110 ( .A(n2410), .ZN(n19891) );
NOR2_X1 U17111 ( .A1(n19912), .A2(n2117), .ZN(n2698) );
NAND2_X1 U17112 ( .A1(n10482), .A2(n10051), .ZN(n10158) );
NOR2_X1 U17113 ( .A1(n19927), .A2(n2117), .ZN(n2455) );
NOR2_X1 U17114 ( .A1(n19934), .A2(n2117), .ZN(n2537) );
INV_X1 U17115 ( .A(n2164), .ZN(n20904) );
INV_X1 U17116 ( .A(n10493), .ZN(n20956) );
NOR2_X1 U17117 ( .A1(n4291), .A2(n20110), .ZN(n4275) );
AND2_X1 U17118 ( .A1(n2554), .A2(n2142), .ZN(n2508) );
NOR2_X1 U17119 ( .A1(n19914), .A2(n2555), .ZN(n2554) );
NOR2_X1 U17120 ( .A1(n2141), .A2(n2556), .ZN(n2555) );
NAND2_X1 U17121 ( .A1(n2410), .A2(n2557), .ZN(n2556) );
NAND2_X1 U17122 ( .A1(n8141), .A2(n5164), .ZN(n7716) );
NOR2_X1 U17123 ( .A1(n7581), .A2(n20988), .ZN(n8141) );
NOR2_X1 U17124 ( .A1(n9837), .A2(n19982), .ZN(n8436) );
INV_X1 U17125 ( .A(n6310), .ZN(n20940) );
NAND2_X1 U17126 ( .A1(n2112), .A2(n2347), .ZN(n2279) );
NAND2_X1 U17127 ( .A1(n2348), .A2(n2349), .ZN(n2347) );
NAND2_X1 U17128 ( .A1(n19906), .A2(n2351), .ZN(n2348) );
NAND2_X1 U17129 ( .A1(n2352), .A2(n19914), .ZN(n2351) );
NAND2_X1 U17130 ( .A1(n19896), .A2(n2112), .ZN(n2590) );
INV_X1 U17131 ( .A(n5088), .ZN(n20992) );
INV_X1 U17132 ( .A(n2349), .ZN(n19897) );
NAND2_X1 U17133 ( .A1(n21305), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N16), .ZN(n21311) );
NOR2_X1 U17134 ( .A1(n21401), .A2(n19870), .ZN(n21305) );
NAND2_X1 U17135 ( .A1(n21312), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N18), .ZN(n21318) );
NOR2_X1 U17136 ( .A1(n21311), .A2(n19865), .ZN(n21312) );
NAND2_X1 U17137 ( .A1(n21319), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N20), .ZN(n21325) );
NOR2_X1 U17138 ( .A1(n21318), .A2(n19860), .ZN(n21319) );
NAND2_X1 U17139 ( .A1(n21326), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N22), .ZN(n21332) );
NOR2_X1 U17140 ( .A1(n21325), .A2(n19855), .ZN(n21326) );
NAND2_X1 U17141 ( .A1(n21333), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N24), .ZN(n21339) );
NOR2_X1 U17142 ( .A1(n21332), .A2(n19850), .ZN(n21333) );
NAND2_X1 U17143 ( .A1(n21340), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N26), .ZN(n21346) );
NOR2_X1 U17144 ( .A1(n21339), .A2(n19845), .ZN(n21340) );
NAND2_X1 U17145 ( .A1(n21347), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N28), .ZN(n21353) );
NOR2_X1 U17146 ( .A1(n21346), .A2(n19840), .ZN(n21347) );
NAND2_X1 U17147 ( .A1(n21354), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N30), .ZN(n21360) );
NOR2_X1 U17148 ( .A1(n21353), .A2(n19835), .ZN(n21354) );
NAND2_X1 U17149 ( .A1(n21361), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N32), .ZN(n21367) );
NOR2_X1 U17150 ( .A1(n21360), .A2(n19830), .ZN(n21361) );
NAND2_X1 U17151 ( .A1(n21368), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N34), .ZN(n21376) );
NOR2_X1 U17152 ( .A1(n21367), .A2(n19825), .ZN(n21368) );
NAND2_X1 U17153 ( .A1(n21304), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N14), .ZN(n21401) );
NOR2_X1 U17154 ( .A1(n21395), .A2(n20725), .ZN(n21304) );
NAND2_X1 U17155 ( .A1(n21303), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N12), .ZN(n21395) );
NOR2_X1 U17156 ( .A1(n21389), .A2(n20736), .ZN(n21303) );
NAND2_X1 U17157 ( .A1(n21302), .A2(n20878), .ZN(n21389) );
NOR2_X1 U17158 ( .A1(n20747), .A2(n16265), .ZN(n21302) );
NAND2_X1 U17159 ( .A1(n10425), .A2(n20932), .ZN(n5138) );
INV_X1 U17160 ( .A(n2112), .ZN(n19941) );
AND2_X1 U17161 ( .A1(n7720), .A2(n19983), .ZN(n7032) );
NAND2_X1 U17162 ( .A1(n1576), .A2(n20993), .ZN(n1541) );
NAND2_X1 U17163 ( .A1(n10051), .A2(n10481), .ZN(n10157) );
NAND2_X1 U17164 ( .A1(n16439), .A2(n1446), .ZN(n3611) );
NOR2_X1 U17165 ( .A1(n16439), .A2(n19853), .ZN(n3526) );
NOR2_X1 U17166 ( .A1(n16439), .A2(n19856), .ZN(n3531) );
NOR2_X1 U17167 ( .A1(n16439), .A2(n19858), .ZN(n3536) );
NOR2_X1 U17168 ( .A1(n16439), .A2(n19861), .ZN(n3541) );
NOR2_X1 U17169 ( .A1(n16439), .A2(n19866), .ZN(n3551) );
NAND2_X1 U17170 ( .A1(n19900), .A2(n2655), .ZN(n2408) );
NAND2_X1 U17171 ( .A1(n2029), .A2(n2655), .ZN(n2384) );
NOR2_X1 U17172 ( .A1(n2024), .A2(n2590), .ZN(n2589) );
NOR2_X1 U17173 ( .A1(n2024), .A2(n2384), .ZN(n2694) );
NAND2_X1 U17174 ( .A1(n10164), .A2(n10165), .ZN(n6235) );
NOR2_X1 U17175 ( .A1(n10170), .A2(n10171), .ZN(n10164) );
NOR2_X1 U17176 ( .A1(n10166), .A2(n10167), .ZN(n10165) );
NOR2_X1 U17177 ( .A1(n10174), .A2(n10175), .ZN(n10170) );
INV_X1 U17178 ( .A(n1395), .ZN(n20945) );
NAND2_X1 U17179 ( .A1(n20985), .A2(n5146), .ZN(n5164) );
NOR2_X1 U17180 ( .A1(n16439), .A2(n3027), .ZN(n3714) );
NAND2_X1 U17181 ( .A1(n19983), .A2(n8074), .ZN(n8079) );
NOR2_X1 U17182 ( .A1(n19931), .A2(n2471), .ZN(n2482) );
NOR2_X1 U17183 ( .A1(n19914), .A2(n2471), .ZN(n2722) );
NOR2_X1 U17184 ( .A1(n16440), .A2(n19838), .ZN(n3485) );
NOR2_X1 U17185 ( .A1(n16441), .A2(n19826), .ZN(n3460) );
NOR2_X1 U17186 ( .A1(n16440), .A2(n19831), .ZN(n3470) );
NOR2_X1 U17187 ( .A1(n16441), .A2(n19833), .ZN(n3475) );
NOR2_X1 U17188 ( .A1(n16440), .A2(n19836), .ZN(n3480) );
NOR2_X1 U17189 ( .A1(n16441), .A2(n19843), .ZN(n3506) );
NOR2_X1 U17190 ( .A1(n16440), .A2(n19846), .ZN(n3511) );
NOR2_X1 U17191 ( .A1(n16439), .A2(n19848), .ZN(n3516) );
NOR2_X1 U17192 ( .A1(n16441), .A2(n20731), .ZN(n3415) );
NOR2_X1 U17193 ( .A1(n16441), .A2(n19813), .ZN(n3430) );
NOR2_X1 U17194 ( .A1(n16441), .A2(n19815), .ZN(n3435) );
NOR2_X1 U17195 ( .A1(n16441), .A2(n19868), .ZN(n3394) );
NOR2_X1 U17196 ( .A1(n16441), .A2(n19871), .ZN(n3400) );
NOR2_X1 U17197 ( .A1(n16441), .A2(n20726), .ZN(n3410) );
NOR2_X1 U17198 ( .A1(n16441), .A2(n20737), .ZN(n3420) );
NOR2_X1 U17199 ( .A1(n16441), .A2(n20720), .ZN(n3405) );
NOR2_X1 U17200 ( .A1(n16440), .A2(n20742), .ZN(n3425) );
NOR2_X1 U17201 ( .A1(n16441), .A2(n20748), .ZN(n3440) );
NOR2_X1 U17202 ( .A1(n16441), .A2(n19818), .ZN(n3445) );
NOR2_X1 U17203 ( .A1(n2725), .A2(n2441), .ZN(n2759) );
NOR2_X1 U17204 ( .A1(n19887), .A2(n2441), .ZN(n2563) );
INV_X1 U17205 ( .A(n2026), .ZN(n19887) );
NOR2_X1 U17206 ( .A1(n2624), .A2(n2409), .ZN(n2629) );
NOR2_X1 U17207 ( .A1(n2015), .A2(n2024), .ZN(n2023) );
NAND2_X1 U17208 ( .A1(n8417), .A2(n19983), .ZN(n8306) );
NOR2_X1 U17209 ( .A1(n8101), .A2(n8312), .ZN(n8417) );
NOR2_X1 U17210 ( .A1(n2152), .A2(n2028), .ZN(n2588) );
INV_X1 U17211 ( .A(n4417), .ZN(n20910) );
NAND2_X1 U17212 ( .A1(n16424), .A2(n4273), .ZN(n4271) );
NOR2_X1 U17213 ( .A1(n10172), .A2(n10175), .ZN(n10207) );
NOR2_X1 U17214 ( .A1(n20757), .A2(n4919), .ZN(n5083) );
NOR2_X1 U17215 ( .A1(n5173), .A2(n5172), .ZN(n5176) );
NOR2_X1 U17216 ( .A1(n19929), .A2(n2638), .ZN(n2628) );
NOR2_X1 U17217 ( .A1(n2332), .A2(n19891), .ZN(n2638) );
NOR2_X1 U17218 ( .A1(n20963), .A2(n10102), .ZN(n10174) );
NOR2_X1 U17219 ( .A1(n2267), .A2(n16454), .ZN(n2264) );
NOR2_X1 U17220 ( .A1(n2268), .A2(n2026), .ZN(n2267) );
AND2_X1 U17221 ( .A1(n2269), .A2(n2270), .ZN(n2268) );
NOR2_X1 U17222 ( .A1(n19927), .A2(n2106), .ZN(n2098) );
NOR2_X1 U17223 ( .A1(n2107), .A2(n2108), .ZN(n2106) );
NAND2_X1 U17224 ( .A1(n2109), .A2(n2110), .ZN(n2108) );
NAND2_X1 U17225 ( .A1(n2111), .A2(n2112), .ZN(n2110) );
NOR2_X1 U17226 ( .A1(n19934), .A2(n2408), .ZN(n2716) );
NOR2_X1 U17227 ( .A1(n19934), .A2(n2202), .ZN(n2219) );
NOR2_X1 U17228 ( .A1(n19931), .A2(n2179), .ZN(n2175) );
NOR2_X1 U17229 ( .A1(n2180), .A2(n2181), .ZN(n2179) );
NAND2_X1 U17230 ( .A1(n2138), .A2(n2036), .ZN(n2181) );
NOR2_X1 U17231 ( .A1(n2406), .A2(n2407), .ZN(n2405) );
NAND2_X1 U17232 ( .A1(n19894), .A2(n2408), .ZN(n2407) );
NAND2_X1 U17233 ( .A1(n2409), .A2(n2410), .ZN(n2406) );
NAND2_X1 U17234 ( .A1(n4425), .A2(n20906), .ZN(n5382) );
NOR2_X1 U17235 ( .A1(n19925), .A2(n2307), .ZN(n2336) );
NOR2_X1 U17236 ( .A1(n19885), .A2(n3567), .ZN(n3578) );
NOR2_X1 U17237 ( .A1(n19923), .A2(n2307), .ZN(n2311) );
NAND2_X1 U17238 ( .A1(n1394), .A2(n1395), .ZN(n1319) );
NOR2_X1 U17239 ( .A1(n2762), .A2(n2763), .ZN(n2761) );
NAND2_X1 U17240 ( .A1(n2768), .A2(n2769), .ZN(n2762) );
NAND2_X1 U17241 ( .A1(n2764), .A2(n2765), .ZN(n2763) );
NAND2_X1 U17242 ( .A1(n19916), .A2(n2770), .ZN(n2769) );
NOR2_X1 U17243 ( .A1(n2484), .A2(n2485), .ZN(n2483) );
NAND2_X1 U17244 ( .A1(n2241), .A2(n2182), .ZN(n2485) );
NOR2_X1 U17245 ( .A1(n19939), .A2(n2349), .ZN(n2484) );
NOR2_X1 U17246 ( .A1(n10199), .A2(n20957), .ZN(n10198) );
INV_X1 U17247 ( .A(n10201), .ZN(n20957) );
NOR2_X1 U17248 ( .A1(n20972), .A2(n10203), .ZN(n10199) );
INV_X1 U17249 ( .A(n10204), .ZN(n20972) );
NOR2_X1 U17250 ( .A1(n2038), .A2(n2039), .ZN(n2037) );
NAND2_X1 U17251 ( .A1(n2044), .A2(n2045), .ZN(n2038) );
NAND2_X1 U17252 ( .A1(n2040), .A2(n2041), .ZN(n2039) );
NAND2_X1 U17253 ( .A1(n2046), .A2(n2047), .ZN(n2045) );
NOR2_X1 U17254 ( .A1(n19984), .A2(n5202), .ZN(n5213) );
NOR2_X1 U17255 ( .A1(n2143), .A2(n16455), .ZN(n2132) );
NOR2_X1 U17256 ( .A1(n2144), .A2(n2145), .ZN(n2143) );
NAND2_X1 U17257 ( .A1(n2146), .A2(n2147), .ZN(n2145) );
NOR2_X1 U17258 ( .A1(n2152), .A2(n19929), .ZN(n2144) );
NOR2_X1 U17259 ( .A1(n2010), .A2(n16454), .ZN(n2006) );
NOR2_X1 U17260 ( .A1(n2011), .A2(n2012), .ZN(n2010) );
NAND2_X1 U17261 ( .A1(n2013), .A2(n2014), .ZN(n2012) );
NOR2_X1 U17262 ( .A1(n19921), .A2(n19902), .ZN(n2011) );
NOR2_X1 U17263 ( .A1(n19780), .A2(n8557), .ZN(n9560) );
INV_X1 U17264 ( .A(n1075), .ZN(n19780) );
NOR2_X1 U17265 ( .A1(n19782), .A2(n16376), .ZN(n9602) );
INV_X1 U17266 ( .A(n1119), .ZN(n19782) );
NOR2_X1 U17267 ( .A1(n19790), .A2(n8557), .ZN(n9754) );
INV_X1 U17268 ( .A(n1275), .ZN(n19790) );
NOR2_X1 U17269 ( .A1(n19810), .A2(n16376), .ZN(n9389) );
INV_X1 U17270 ( .A(n904), .ZN(n19810) );
NAND2_X1 U17271 ( .A1(n16448), .A2(n2164), .ZN(n2755) );
NAND2_X1 U17272 ( .A1(n16422), .A2(n4273), .ZN(n4279) );
INV_X1 U17273 ( .A(n1565), .ZN(n20935) );
NOR2_X1 U17274 ( .A1(n19804), .A2(n8557), .ZN(n8780) );
INV_X1 U17275 ( .A(n301), .ZN(n19804) );
NOR2_X1 U17276 ( .A1(n19806), .A2(n8557), .ZN(n8826) );
INV_X1 U17277 ( .A(n342), .ZN(n19806) );
NOR2_X1 U17278 ( .A1(n19752), .A2(n8557), .ZN(n8929) );
INV_X1 U17279 ( .A(n427), .ZN(n19752) );
NOR2_X1 U17280 ( .A1(n19802), .A2(n8557), .ZN(n8736) );
INV_X1 U17281 ( .A(n260), .ZN(n19802) );
NAND2_X1 U17282 ( .A1(n1561), .A2(n1562), .ZN(n1544) );
OR2_X1 U17283 ( .A1(n16463), .A2(n1564), .ZN(n1562) );
NAND2_X1 U17284 ( .A1(n1565), .A2(n1566), .ZN(n1561) );
INV_X1 U17285 ( .A(n5120), .ZN(n20989) );
NAND2_X1 U17286 ( .A1(n21377), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N36), .ZN(n21380) );
NOR2_X1 U17287 ( .A1(n21376), .A2(n19820), .ZN(n21377) );
NAND2_X1 U17288 ( .A1(n4260), .A2(n20906), .ZN(n4067) );
NOR2_X1 U17289 ( .A1(n4258), .A2(n20763), .ZN(n4260) );
NAND2_X1 U17290 ( .A1(n4256), .A2(n20906), .ZN(n4066) );
NOR2_X1 U17291 ( .A1(n4257), .A2(n4258), .ZN(n4256) );
NAND2_X1 U17292 ( .A1(n2714), .A2(n19919), .ZN(n2666) );
NOR2_X1 U17293 ( .A1(n19917), .A2(n2715), .ZN(n2714) );
NOR2_X1 U17294 ( .A1(n7581), .A2(n7582), .ZN(n7578) );
NOR2_X1 U17295 ( .A1(n19749), .A2(n7562), .ZN(n7582) );
NOR2_X1 U17296 ( .A1(n5169), .A2(n5170), .ZN(n5165) );
NOR2_X1 U17297 ( .A1(n20930), .A2(n5172), .ZN(n5170) );
INV_X1 U17298 ( .A(n5173), .ZN(n20930) );
NOR2_X1 U17299 ( .A1(n4020), .A2(n7589), .ZN(n7587) );
NOR2_X1 U17300 ( .A1(n19803), .A2(n7562), .ZN(n7589) );
NOR2_X1 U17301 ( .A1(n2621), .A2(n2622), .ZN(n2615) );
NOR2_X1 U17302 ( .A1(n19934), .A2(n2590), .ZN(n2622) );
NOR2_X1 U17303 ( .A1(n19901), .A2(n2624), .ZN(n2621) );
INV_X1 U17304 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N9), .ZN(n20747) );
INV_X1 U17305 ( .A(n5249), .ZN(n20932) );
NAND2_X1 U17306 ( .A1(n5085), .A2(n4417), .ZN(n4936) );
AND2_X1 U17307 ( .A1(n1420), .A2(n1423), .ZN(n5085) );
INV_X1 U17308 ( .A(n1597), .ZN(n20938) );
NAND2_X1 U17309 ( .A1(n2773), .A2(n19914), .ZN(n2523) );
INV_X1 U17310 ( .A(n5096), .ZN(n21001) );
INV_X1 U17311 ( .A(n1687), .ZN(n20994) );
NAND2_X1 U17312 ( .A1(n4955), .A2(n4417), .ZN(n4797) );
AND2_X1 U17313 ( .A1(n1423), .A2(n1422), .ZN(n4955) );
NAND2_X1 U17314 ( .A1(n10505), .A2(n10156), .ZN(n10060) );
NAND2_X1 U17315 ( .A1(n19897), .A2(n2112), .ZN(n2235) );
NAND2_X1 U17316 ( .A1(n19897), .A2(n2270), .ZN(n2582) );
NAND2_X1 U17317 ( .A1(n2182), .A2(n2183), .ZN(n2059) );
NAND2_X1 U17318 ( .A1(n2112), .A2(n2184), .ZN(n2183) );
NAND2_X1 U17319 ( .A1(n19923), .A2(n2720), .ZN(n2048) );
NAND2_X1 U17320 ( .A1(n8415), .A2(n8416), .ZN(n8414) );
NAND2_X1 U17321 ( .A1(n8310), .A2(n19980), .ZN(n8416) );
NAND2_X1 U17322 ( .A1(n8313), .A2(n8306), .ZN(n8415) );
AND2_X1 U17323 ( .A1(n4417), .A2(n4418), .ZN(n4410) );
NAND2_X1 U17324 ( .A1(n20908), .A2(n4420), .ZN(n4418) );
NAND2_X1 U17325 ( .A1(n4421), .A2(n4422), .ZN(n4420) );
INV_X1 U17326 ( .A(n4412), .ZN(n20908) );
NAND2_X1 U17327 ( .A1(n2270), .A2(n2269), .ZN(n2346) );
INV_X1 U17328 ( .A(n1416), .ZN(n20937) );
NAND2_X1 U17329 ( .A1(n19890), .A2(n2270), .ZN(n2147) );
NAND2_X1 U17330 ( .A1(n19906), .A2(n2388), .ZN(n2356) );
NAND2_X1 U17331 ( .A1(n10512), .A2(n20956), .ZN(n10504) );
NOR2_X1 U17332 ( .A1(n10156), .A2(n10501), .ZN(n10512) );
NAND2_X1 U17333 ( .A1(n10161), .A2(n20942), .ZN(n10127) );
NOR2_X1 U17334 ( .A1(n20944), .A2(n6306), .ZN(n10161) );
INV_X1 U17335 ( .A(n5735), .ZN(n20921) );
NAND2_X1 U17336 ( .A1(n20936), .A2(n8557), .ZN(n9973) );
NAND2_X1 U17337 ( .A1(n7081), .A2(n7082), .ZN(n7072) );
NOR2_X1 U17338 ( .A1(n16201), .A2(n7084), .ZN(n7081) );
INV_X1 U17339 ( .A(n3126), .ZN(n19873) );
NAND2_X1 U17340 ( .A1(n4916), .A2(n16424), .ZN(n4915) );
NAND2_X1 U17341 ( .A1(n4897), .A2(n16424), .ZN(n4896) );
NAND2_X1 U17342 ( .A1(n4878), .A2(n16424), .ZN(n4877) );
NAND2_X1 U17343 ( .A1(n4859), .A2(n16424), .ZN(n4858) );
NAND2_X1 U17344 ( .A1(n4840), .A2(n16424), .ZN(n4839) );
NAND2_X1 U17345 ( .A1(n4821), .A2(n16424), .ZN(n4820) );
AND2_X1 U17346 ( .A1(n6699), .A2(n4005), .ZN(n3740) );
NOR2_X1 U17347 ( .A1(n6701), .A2(n4046), .ZN(n6699) );
AND2_X1 U17348 ( .A1(n10191), .A2(n20963), .ZN(n10095) );
NOR2_X1 U17349 ( .A1(n10192), .A2(n10193), .ZN(n10191) );
NOR2_X1 U17350 ( .A1(n20973), .A2(n20974), .ZN(n10192) );
AND2_X1 U17351 ( .A1(n2687), .A2(n19917), .ZN(n2139) );
NOR2_X1 U17352 ( .A1(n16457), .A2(n19902), .ZN(n2687) );
AND2_X1 U17353 ( .A1(n2235), .A2(n2850), .ZN(n2725) );
NAND2_X1 U17354 ( .A1(n19917), .A2(n2055), .ZN(n2850) );
AND2_X1 U17355 ( .A1(n7033), .A2(n8106), .ZN(n7795) );
AND2_X1 U17356 ( .A1(n6232), .A2(n6233), .ZN(n1394) );
NOR2_X1 U17357 ( .A1(n6234), .A2(n6235), .ZN(n6232) );
NOR2_X1 U17358 ( .A1(n20952), .A2(n20940), .ZN(n6233) );
NAND2_X1 U17359 ( .A1(n19982), .A2(n8452), .ZN(n8456) );
NAND2_X1 U17360 ( .A1(n5529), .A2(n4425), .ZN(n5385) );
NOR2_X1 U17361 ( .A1(n20085), .A2(n5374), .ZN(n5529) );
NAND2_X1 U17362 ( .A1(n20988), .A2(n20880), .ZN(n7876) );
INV_X1 U17363 ( .A(n4940), .ZN(n20919) );
NAND2_X1 U17364 ( .A1(n8078), .A2(n7041), .ZN(n10317) );
NAND2_X1 U17365 ( .A1(n7023), .A2(n7031), .ZN(n6719) );
NAND2_X1 U17366 ( .A1(n7032), .A2(n7033), .ZN(n7031) );
INV_X1 U17367 ( .A(n10156), .ZN(n20964) );
NAND2_X1 U17368 ( .A1(n4395), .A2(n16422), .ZN(n4399) );
NAND2_X1 U17369 ( .A1(n4376), .A2(n16422), .ZN(n4380) );
NAND2_X1 U17370 ( .A1(n4357), .A2(n16422), .ZN(n4361) );
NAND2_X1 U17371 ( .A1(n4338), .A2(n16422), .ZN(n4342) );
NAND2_X1 U17372 ( .A1(n4319), .A2(n16422), .ZN(n4323) );
NAND2_X1 U17373 ( .A1(n4300), .A2(n16422), .ZN(n4304) );
NAND2_X1 U17374 ( .A1(n2053), .A2(n2054), .ZN(n2030) );
NOR2_X1 U17375 ( .A1(n2059), .A2(n2060), .ZN(n2053) );
NOR2_X1 U17376 ( .A1(n2055), .A2(n2056), .ZN(n2054) );
NOR2_X1 U17377 ( .A1(n19894), .A2(n2058), .ZN(n2056) );
NAND2_X1 U17378 ( .A1(n5224), .A2(n5225), .ZN(n2003) );
NOR2_X1 U17379 ( .A1(n5226), .A2(n5141), .ZN(n5224) );
NOR2_X1 U17380 ( .A1(n5184), .A2(n5222), .ZN(n5226) );
NAND2_X1 U17381 ( .A1(n3054), .A2(n3055), .ZN(n3041) );
NAND2_X1 U17382 ( .A1(n1447), .A2(n16439), .ZN(n3055) );
AND2_X1 U17383 ( .A1(n2395), .A2(n2396), .ZN(n2383) );
NOR2_X1 U17384 ( .A1(n2400), .A2(n2401), .ZN(n2395) );
NOR2_X1 U17385 ( .A1(n2397), .A2(n2398), .ZN(n2396) );
NOR2_X1 U17386 ( .A1(n19912), .A2(n19940), .ZN(n2401) );
NAND2_X1 U17387 ( .A1(n2700), .A2(n2701), .ZN(n2682) );
AND2_X1 U17388 ( .A1(n2303), .A2(n2666), .ZN(n2700) );
NAND2_X1 U17389 ( .A1(n2702), .A2(n19905), .ZN(n2701) );
AND2_X1 U17390 ( .A1(n2668), .A2(n2669), .ZN(n2242) );
NOR2_X1 U17391 ( .A1(n2670), .A2(n2671), .ZN(n2668) );
NOR2_X1 U17392 ( .A1(n19942), .A2(n16456), .ZN(n2671) );
NOR2_X1 U17393 ( .A1(n2673), .A2(n19881), .ZN(n2670) );
AND2_X1 U17394 ( .A1(n2494), .A2(n2495), .ZN(n2071) );
NAND2_X1 U17395 ( .A1(n19875), .A2(n2496), .ZN(n2495) );
NOR2_X1 U17396 ( .A1(n2339), .A2(n2508), .ZN(n2494) );
NAND2_X1 U17397 ( .A1(n2497), .A2(n2498), .ZN(n2496) );
AND2_X1 U17398 ( .A1(n2460), .A2(n2461), .ZN(n2064) );
NOR2_X1 U17399 ( .A1(n2462), .A2(n2463), .ZN(n2460) );
NOR2_X1 U17400 ( .A1(n19929), .A2(n2471), .ZN(n2462) );
NOR2_X1 U17401 ( .A1(n2464), .A2(n19881), .ZN(n2463) );
AND2_X1 U17402 ( .A1(n2451), .A2(n2452), .ZN(n2061) );
NOR2_X1 U17403 ( .A1(n2454), .A2(n2455), .ZN(n2451) );
NAND2_X1 U17404 ( .A1(n2142), .A2(n2453), .ZN(n2452) );
NOR2_X1 U17405 ( .A1(n2456), .A2(n2457), .ZN(n2454) );
AND2_X1 U17406 ( .A1(n2612), .A2(n2613), .ZN(n2090) );
NAND2_X1 U17407 ( .A1(n16452), .A2(n2614), .ZN(n2613) );
NAND2_X1 U17408 ( .A1(n2142), .A2(n2625), .ZN(n2612) );
NAND2_X1 U17409 ( .A1(n2615), .A2(n2616), .ZN(n2614) );
AND2_X1 U17410 ( .A1(n2669), .A2(n2448), .ZN(n2412) );
NAND2_X1 U17411 ( .A1(n2387), .A2(n2055), .ZN(n2266) );
AND2_X1 U17412 ( .A1(n2388), .A2(n16453), .ZN(n2387) );
AND2_X1 U17413 ( .A1(n16423), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_11), .ZN(n4891) );
AND2_X1 U17414 ( .A1(n16423), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_12), .ZN(n4872) );
AND2_X1 U17415 ( .A1(n4275), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_14), .ZN(n4834) );
AND2_X1 U17416 ( .A1(n16423), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_9), .ZN(n4264) );
INV_X1 U17417 ( .A(n4257), .ZN(n20763) );
INV_X1 U17418 ( .A(n4431), .ZN(n21003) );
NAND2_X1 U17419 ( .A1(n20949), .A2(n10134), .ZN(n8601) );
INV_X1 U17420 ( .A(n4258), .ZN(n20999) );
INV_X1 U17421 ( .A(n10051), .ZN(n20950) );
NAND2_X1 U17422 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N37), .A2(n19817), .ZN(n21381) );
INV_X1 U17423 ( .A(n21380), .ZN(n19817) );
NAND2_X1 U17424 ( .A1(n4449), .A2(n4272), .ZN(n4448) );
NAND2_X1 U17425 ( .A1(n4802), .A2(n4272), .ZN(n4801) );
NAND2_X1 U17426 ( .A1(n4780), .A2(n16424), .ZN(n4779) );
NAND2_X1 U17427 ( .A1(n4759), .A2(n4272), .ZN(n4758) );
NAND2_X1 U17428 ( .A1(n4738), .A2(n16424), .ZN(n4737) );
NAND2_X1 U17429 ( .A1(n4699), .A2(n4272), .ZN(n4698) );
NAND2_X1 U17430 ( .A1(n4678), .A2(n16424), .ZN(n4677) );
NAND2_X1 U17431 ( .A1(n4657), .A2(n4272), .ZN(n4656) );
NAND2_X1 U17432 ( .A1(n4636), .A2(n16424), .ZN(n4635) );
NAND2_X1 U17433 ( .A1(n4615), .A2(n4272), .ZN(n4614) );
NAND2_X1 U17434 ( .A1(n4594), .A2(n16424), .ZN(n4593) );
NAND2_X1 U17435 ( .A1(n4573), .A2(n4272), .ZN(n4572) );
NAND2_X1 U17436 ( .A1(n4552), .A2(n4272), .ZN(n4551) );
NAND2_X1 U17437 ( .A1(n4531), .A2(n4272), .ZN(n4530) );
NAND2_X1 U17438 ( .A1(n4510), .A2(n4272), .ZN(n4509) );
NAND2_X1 U17439 ( .A1(n4470), .A2(n4272), .ZN(n4469) );
NAND2_X1 U17440 ( .A1(n4718), .A2(n16424), .ZN(n4717) );
NAND2_X1 U17441 ( .A1(n4489), .A2(n4272), .ZN(n4488) );
NAND2_X1 U17442 ( .A1(n4395), .A2(n4272), .ZN(n4394) );
NAND2_X1 U17443 ( .A1(n4376), .A2(n16424), .ZN(n4375) );
NAND2_X1 U17444 ( .A1(n4357), .A2(n4272), .ZN(n4356) );
NAND2_X1 U17445 ( .A1(n4338), .A2(n16424), .ZN(n4337) );
NAND2_X1 U17446 ( .A1(n4319), .A2(n4272), .ZN(n4318) );
NAND2_X1 U17447 ( .A1(n4300), .A2(n16424), .ZN(n4299) );
NAND2_X1 U17448 ( .A1(n4916), .A2(n4280), .ZN(n4923) );
NAND2_X1 U17449 ( .A1(n4449), .A2(n4280), .ZN(n4453) );
NAND2_X1 U17450 ( .A1(n4897), .A2(n16422), .ZN(n4901) );
NAND2_X1 U17451 ( .A1(n4878), .A2(n4280), .ZN(n4882) );
NAND2_X1 U17452 ( .A1(n4859), .A2(n16422), .ZN(n4863) );
NAND2_X1 U17453 ( .A1(n4840), .A2(n4280), .ZN(n4844) );
NAND2_X1 U17454 ( .A1(n4821), .A2(n16422), .ZN(n4825) );
NAND2_X1 U17455 ( .A1(n4802), .A2(n4280), .ZN(n4806) );
NAND2_X1 U17456 ( .A1(n4780), .A2(n16422), .ZN(n4784) );
NAND2_X1 U17457 ( .A1(n4759), .A2(n4280), .ZN(n4763) );
NAND2_X1 U17458 ( .A1(n4738), .A2(n16422), .ZN(n4742) );
NAND2_X1 U17459 ( .A1(n4699), .A2(n4280), .ZN(n4703) );
NAND2_X1 U17460 ( .A1(n4678), .A2(n4280), .ZN(n4682) );
NAND2_X1 U17461 ( .A1(n4657), .A2(n4280), .ZN(n4661) );
NAND2_X1 U17462 ( .A1(n4636), .A2(n4280), .ZN(n4640) );
NAND2_X1 U17463 ( .A1(n4615), .A2(n4280), .ZN(n4619) );
NAND2_X1 U17464 ( .A1(n4594), .A2(n4280), .ZN(n4598) );
NAND2_X1 U17465 ( .A1(n4573), .A2(n16422), .ZN(n4577) );
NAND2_X1 U17466 ( .A1(n4552), .A2(n4280), .ZN(n4556) );
NAND2_X1 U17467 ( .A1(n4531), .A2(n16422), .ZN(n4535) );
NAND2_X1 U17468 ( .A1(n4510), .A2(n4280), .ZN(n4514) );
NAND2_X1 U17469 ( .A1(n4470), .A2(n16422), .ZN(n4474) );
NAND2_X1 U17470 ( .A1(n4718), .A2(n16422), .ZN(n4722) );
NAND2_X1 U17471 ( .A1(n4489), .A2(n4280), .ZN(n4493) );
INV_X1 U17472 ( .A(n7580), .ZN(n20924) );
INV_X1 U17473 ( .A(n5222), .ZN(n19985) );
INV_X1 U17474 ( .A(n2522), .ZN(n19909) );
INV_X1 U17475 ( .A(n5210), .ZN(n19984) );
INV_X1 U17476 ( .A(n1446), .ZN(n20878) );
NAND2_X1 U17477 ( .A1(n7032), .A2(n7571), .ZN(n7570) );
NAND2_X1 U17478 ( .A1(n1411), .A2(n6230), .ZN(n5826) );
NAND2_X1 U17479 ( .A1(n1342), .A2(n6231), .ZN(n6230) );
AND2_X1 U17480 ( .A1(n4425), .A2(n5091), .ZN(n5818) );
INV_X1 U17481 ( .A(n5091), .ZN(n20961) );
NAND2_X1 U17482 ( .A1(n5378), .A2(n21004), .ZN(n5278) );
NOR2_X1 U17483 ( .A1(n21003), .A2(n5374), .ZN(n5378) );
NAND2_X1 U17484 ( .A1(n2539), .A2(n2029), .ZN(n2765) );
INV_X1 U17485 ( .A(n6234), .ZN(n20943) );
INV_X1 U17486 ( .A(n2060), .ZN(n19901) );
AND2_X1 U17487 ( .A1(n4924), .A2(n16424), .ZN(n4280) );
NOR2_X1 U17488 ( .A1(n21002), .A2(n20910), .ZN(n4924) );
INV_X1 U17489 ( .A(n10234), .ZN(n20965) );
INV_X1 U17490 ( .A(n2697), .ZN(n19896) );
INV_X1 U17491 ( .A(n10134), .ZN(n20948) );
INV_X1 U17492 ( .A(n5571), .ZN(n20911) );
INV_X1 U17493 ( .A(n10330), .ZN(n20933) );
NAND2_X1 U17494 ( .A1(n20943), .A2(n6306), .ZN(n10089) );
INV_X1 U17495 ( .A(n5153), .ZN(n20873) );
NAND2_X1 U17496 ( .A1(n2666), .A2(n2303), .ZN(n2712) );
NAND2_X1 U17497 ( .A1(n6231), .A2(n1395), .ZN(n10118) );
INV_X1 U17498 ( .A(n5716), .ZN(n20922) );
INV_X1 U17499 ( .A(n5267), .ZN(n20936) );
NAND2_X1 U17500 ( .A1(n2182), .A2(n2399), .ZN(n2398) );
INV_X1 U17501 ( .A(n7705), .ZN(n20915) );
AND2_X1 U17502 ( .A1(n8452), .A2(n8883), .ZN(n8455) );
AND2_X1 U17503 ( .A1(n5372), .A2(n21003), .ZN(n5277) );
NOR2_X1 U17504 ( .A1(n20110), .A2(n5374), .ZN(n5372) );
NAND2_X1 U17505 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N9), .A2(n1446), .ZN(n21375) );
NAND2_X1 U17506 ( .A1(n8308), .A2(n8309), .ZN(n8165) );
OR2_X1 U17507 ( .A1(n8313), .A2(n19980), .ZN(n8308) );
NAND2_X1 U17508 ( .A1(n8310), .A2(n20851), .ZN(n8309) );
INV_X1 U17509 ( .A(n8312), .ZN(n20851) );
NAND2_X1 U17510 ( .A1(n2686), .A2(n2702), .ZN(n2719) );
NAND2_X1 U17511 ( .A1(n8111), .A2(n8112), .ZN(n8107) );
NAND2_X1 U17512 ( .A1(n8113), .A2(n20853), .ZN(n8112) );
NOR2_X1 U17513 ( .A1(n7720), .A2(n8116), .ZN(n8111) );
NAND2_X1 U17514 ( .A1(n20868), .A2(n8115), .ZN(n8113) );
NAND2_X1 U17515 ( .A1(n20973), .A2(n20963), .ZN(n10213) );
NAND2_X1 U17516 ( .A1(n2177), .A2(n19879), .ZN(n2176) );
OR2_X1 U17517 ( .A1(n2104), .A2(n19927), .ZN(n2177) );
NAND2_X1 U17518 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N13), .A2(n21395), .ZN(n21393) );
NAND2_X1 U17519 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N15), .A2(n21401), .ZN(n21399) );
NAND2_X1 U17520 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N17), .A2(n21311), .ZN(n21306) );
NAND2_X1 U17521 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N19), .A2(n21318), .ZN(n21313) );
NAND2_X1 U17522 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N21), .A2(n21325), .ZN(n21320) );
NAND2_X1 U17523 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N23), .A2(n21332), .ZN(n21327) );
NAND2_X1 U17524 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N25), .A2(n21339), .ZN(n21334) );
NAND2_X1 U17525 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N27), .A2(n21346), .ZN(n21341) );
NAND2_X1 U17526 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N29), .A2(n21353), .ZN(n21348) );
NAND2_X1 U17527 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N31), .A2(n21360), .ZN(n21355) );
NAND2_X1 U17528 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N33), .A2(n21367), .ZN(n21362) );
NAND2_X1 U17529 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N35), .A2(n21376), .ZN(n21369) );
NAND2_X1 U17530 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N11), .A2(n21389), .ZN(n21387) );
NAND2_X1 U17531 ( .A1(n2313), .A2(n19880), .ZN(n2312) );
NAND2_X1 U17532 ( .A1(n16451), .A2(n2315), .ZN(n2313) );
NAND2_X1 U17533 ( .A1(n2316), .A2(n2152), .ZN(n2315) );
NOR2_X1 U17534 ( .A1(n19895), .A2(n2318), .ZN(n2316) );
NAND2_X1 U17535 ( .A1(n2338), .A2(n19880), .ZN(n2337) );
NAND2_X1 U17536 ( .A1(n2340), .A2(n19899), .ZN(n2338) );
NOR2_X1 U17537 ( .A1(n19929), .A2(n19881), .ZN(n2340) );
INV_X1 U17538 ( .A(n4919), .ZN(n20023) );
NAND2_X1 U17539 ( .A1(n2771), .A2(n2772), .ZN(n2770) );
NAND2_X1 U17540 ( .A1(n2539), .A2(n2049), .ZN(n2772) );
NOR2_X1 U17541 ( .A1(n19895), .A2(n2797), .ZN(n2771) );
NOR2_X1 U17542 ( .A1(n2523), .A2(n2582), .ZN(n2797) );
NAND2_X1 U17543 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N37), .A2(n21380), .ZN(n21378) );
INV_X1 U17544 ( .A(n5250), .ZN(n20968) );
INV_X1 U17545 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N15), .ZN(n19870) );
INV_X1 U17546 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N17), .ZN(n19865) );
INV_X1 U17547 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N19), .ZN(n19860) );
INV_X1 U17548 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N21), .ZN(n19855) );
INV_X1 U17549 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N25), .ZN(n19845) );
INV_X1 U17550 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N27), .ZN(n19840) );
INV_X1 U17551 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N29), .ZN(n19835) );
INV_X1 U17552 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N31), .ZN(n19830) );
INV_X1 U17553 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N33), .ZN(n19825) );
INV_X1 U17554 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N35), .ZN(n19820) );
INV_X1 U17555 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N11), .ZN(n20736) );
INV_X1 U17556 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N13), .ZN(n20725) );
NAND2_X1 U17557 ( .A1(n5169), .A2(n5198), .ZN(n5191) );
INV_X1 U17558 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N23), .ZN(n19850) );
INV_X1 U17559 ( .A(n6701), .ZN(n20931) );
NAND2_X1 U17560 ( .A1(n20973), .A2(n10256), .ZN(n10255) );
NAND2_X1 U17561 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N12), .A2(n21390), .ZN(n21391) );
NAND2_X1 U17562 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N14), .A2(n21396), .ZN(n21397) );
NAND2_X1 U17563 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N16), .A2(n21402), .ZN(n21403) );
NAND2_X1 U17564 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N18), .A2(n21308), .ZN(n21309) );
NAND2_X1 U17565 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N20), .A2(n21315), .ZN(n21316) );
NAND2_X1 U17566 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N22), .A2(n21322), .ZN(n21323) );
NAND2_X1 U17567 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N24), .A2(n21329), .ZN(n21330) );
NAND2_X1 U17568 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N26), .A2(n21336), .ZN(n21337) );
NAND2_X1 U17569 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N28), .A2(n21343), .ZN(n21344) );
NAND2_X1 U17570 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N30), .A2(n21350), .ZN(n21351) );
NAND2_X1 U17571 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N32), .A2(n21357), .ZN(n21358) );
NAND2_X1 U17572 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N34), .A2(n21364), .ZN(n21365) );
NAND2_X1 U17573 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N36), .A2(n21371), .ZN(n21372) );
NAND2_X1 U17574 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N38), .A2(n21381), .ZN(n21382) );
NAND2_X1 U17575 ( .A1(n20984), .A2(n5216), .ZN(n5215) );
NAND2_X1 U17576 ( .A1(n5198), .A2(n5202), .ZN(n5216) );
NAND2_X1 U17577 ( .A1(n2710), .A2(n2711), .ZN(n2709) );
NOR2_X1 U17578 ( .A1(n2716), .A2(n2717), .ZN(n2710) );
NOR2_X1 U17579 ( .A1(n19904), .A2(n2712), .ZN(n2711) );
NAND2_X1 U17580 ( .A1(n2718), .A2(n2719), .ZN(n2717) );
NAND2_X1 U17581 ( .A1(n2514), .A2(n2515), .ZN(n2513) );
NOR2_X1 U17582 ( .A1(n2520), .A2(n2521), .ZN(n2514) );
NOR2_X1 U17583 ( .A1(n2516), .A2(n2517), .ZN(n2515) );
NOR2_X1 U17584 ( .A1(n19923), .A2(n2522), .ZN(n2521) );
NAND2_X1 U17585 ( .A1(n2626), .A2(n2627), .ZN(n2625) );
NOR2_X1 U17586 ( .A1(n2639), .A2(n2566), .ZN(n2626) );
NOR2_X1 U17587 ( .A1(n2628), .A2(n2629), .ZN(n2627) );
NOR2_X1 U17588 ( .A1(n19925), .A2(n2522), .ZN(n2639) );
NAND2_X1 U17589 ( .A1(n2477), .A2(n19893), .ZN(n2476) );
INV_X1 U17590 ( .A(n2238), .ZN(n19893) );
NOR2_X1 U17591 ( .A1(n19900), .A2(n2480), .ZN(n2477) );
NOR2_X1 U17592 ( .A1(n19931), .A2(n2409), .ZN(n2480) );
NAND2_X1 U17593 ( .A1(n2148), .A2(n19896), .ZN(n2146) );
NOR2_X1 U17594 ( .A1(n19919), .A2(n19940), .ZN(n2148) );
NAND2_X1 U17595 ( .A1(n21384), .A2(n16265), .ZN(n21386) );
AND2_X1 U17596 ( .A1(n16423), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_10), .ZN(n4910) );
AND2_X1 U17597 ( .A1(n4275), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_13), .ZN(n4853) );
AND2_X1 U17598 ( .A1(n4275), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_15), .ZN(n4815) );
AND2_X1 U17599 ( .A1(n16423), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_1), .ZN(n4712) );
AND2_X1 U17600 ( .A1(n16423), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_2), .ZN(n4483) );
AND2_X1 U17601 ( .A1(n4275), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_3), .ZN(n4389) );
AND2_X1 U17602 ( .A1(n16423), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_4), .ZN(n4370) );
AND2_X1 U17603 ( .A1(n16423), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_5), .ZN(n4351) );
AND2_X1 U17604 ( .A1(n16423), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_6), .ZN(n4332) );
AND2_X1 U17605 ( .A1(n16423), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_7), .ZN(n4313) );
OR2_X1 U17606 ( .A1(n16252), .A2(n10108), .ZN(n10160) );
OR2_X1 U17607 ( .A1(n1395), .A2(n6231), .ZN(n16252) );
OR2_X1 U17608 ( .A1(n21389), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N11), .ZN(n21388) );
OR2_X1 U17609 ( .A1(n21395), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N13), .ZN(n21394) );
OR2_X1 U17610 ( .A1(n21401), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N15), .ZN(n21400) );
OR2_X1 U17611 ( .A1(n21311), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N17), .ZN(n21307) );
OR2_X1 U17612 ( .A1(n21318), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N19), .ZN(n21314) );
OR2_X1 U17613 ( .A1(n21325), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N21), .ZN(n21321) );
OR2_X1 U17614 ( .A1(n21332), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N23), .ZN(n21328) );
OR2_X1 U17615 ( .A1(n21339), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N25), .ZN(n21335) );
OR2_X1 U17616 ( .A1(n21346), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N27), .ZN(n21342) );
OR2_X1 U17617 ( .A1(n21353), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N29), .ZN(n21349) );
OR2_X1 U17618 ( .A1(n21360), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N31), .ZN(n21356) );
OR2_X1 U17619 ( .A1(n21367), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N33), .ZN(n21363) );
OR2_X1 U17620 ( .A1(n21376), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N35), .ZN(n21370) );
OR2_X1 U17621 ( .A1(n21380), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N37), .ZN(n21379) );
OR2_X1 U17622 ( .A1(n21390), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N12), .ZN(n21392) );
OR2_X1 U17623 ( .A1(n21396), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N14), .ZN(n21398) );
OR2_X1 U17624 ( .A1(n21402), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N16), .ZN(n21404) );
OR2_X1 U17625 ( .A1(n21308), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N18), .ZN(n21310) );
OR2_X1 U17626 ( .A1(n21315), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N20), .ZN(n21317) );
OR2_X1 U17627 ( .A1(n21322), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N22), .ZN(n21324) );
OR2_X1 U17628 ( .A1(n21329), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N24), .ZN(n21331) );
OR2_X1 U17629 ( .A1(n21336), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N26), .ZN(n21338) );
OR2_X1 U17630 ( .A1(n21343), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N28), .ZN(n21345) );
OR2_X1 U17631 ( .A1(n21350), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N30), .ZN(n21352) );
OR2_X1 U17632 ( .A1(n21357), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N32), .ZN(n21359) );
OR2_X1 U17633 ( .A1(n21364), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N34), .ZN(n21366) );
OR2_X1 U17634 ( .A1(n21371), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N36), .ZN(n21373) );
OR2_X1 U17635 ( .A1(n21381), .A2(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N38), .ZN(n21383) );
OR2_X1 U17636 ( .A1(n2015), .A2(n19931), .ZN(n2014) );
OR2_X1 U17637 ( .A1(n16265), .A2(n21384), .ZN(n21385) );
INV_X1 U17638 ( .A(n2566), .ZN(n19892) );
NOR2_X1 U17639 ( .A1(n5153), .A2(n5154), .ZN(n15555) );
NOR2_X1 U17640 ( .A1(n5155), .A2(n5156), .ZN(n5154) );
NAND2_X1 U17641 ( .A1(n5157), .A2(n19968), .ZN(n5156) );
NAND2_X1 U17642 ( .A1(n5165), .A2(n5166), .ZN(n5155) );
INV_X1 U17643 ( .A(n9837), .ZN(n19981) );
OR2_X1 U17644 ( .A1(n16445), .A2(n16459), .ZN(n2900) );
OR2_X1 U17645 ( .A1(n16445), .A2(n1708), .ZN(n2901) );
INV_X1 U17646 ( .A(n590), .ZN(n19758) );
INV_X1 U17647 ( .A(n630), .ZN(n19760) );
INV_X1 U17648 ( .A(n669), .ZN(n19762) );
INV_X1 U17649 ( .A(n707), .ZN(n19764) );
INV_X1 U17650 ( .A(n744), .ZN(n19766) );
INV_X1 U17651 ( .A(n782), .ZN(n19768) );
INV_X1 U17652 ( .A(n859), .ZN(n19772) );
INV_X1 U17653 ( .A(n940), .ZN(n19774) );
INV_X1 U17654 ( .A(n979), .ZN(n19776) );
INV_X1 U17655 ( .A(n1158), .ZN(n19784) );
INV_X1 U17656 ( .A(n1197), .ZN(n19786) );
INV_X1 U17657 ( .A(n1236), .ZN(n19788) );
INV_X1 U17658 ( .A(n1331), .ZN(n19792) );
INV_X1 U17659 ( .A(n79), .ZN(n19794) );
INV_X1 U17660 ( .A(n127), .ZN(n19796) );
INV_X1 U17661 ( .A(n218), .ZN(n19800) );
INV_X1 U17662 ( .A(n175), .ZN(n19798) );
INV_X1 U17663 ( .A(n1415), .ZN(n19812) );
INV_X1 U17664 ( .A(n472), .ZN(n19808) );
INV_X1 U17665 ( .A(n550), .ZN(n19756) );
INV_X1 U17666 ( .A(n510), .ZN(n19754) );
INV_X1 U17667 ( .A(n383), .ZN(n19750) );
INV_X1 U17668 ( .A(n820), .ZN(n19770) );
INV_X1 U17669 ( .A(n1017), .ZN(n19778) );
INV_X1 U17670 ( .A(n5159), .ZN(n19968) );
NAND2_X1 U17671 ( .A1(n2290), .A2(n2291), .ZN(n15594) );
NOR2_X1 U17672 ( .A1(n2304), .A2(n2305), .ZN(n2290) );
NOR2_X1 U17673 ( .A1(n19877), .A2(n2292), .ZN(n2291) );
NOR2_X1 U17674 ( .A1(n19921), .A2(n2307), .ZN(n2304) );
NAND2_X1 U17675 ( .A1(n6505), .A2(n6506), .ZN(data_req_o) );
NOR2_X1 U17676 ( .A1(n20996), .A2(n6508), .ZN(n6505) );
NOR2_X1 U17677 ( .A1(n20998), .A2(n20995), .ZN(n6506) );
AND2_X1 U17678 ( .A1(n1579), .A2(n1576), .ZN(n6508) );
NAND2_X1 U17679 ( .A1(n2262), .A2(n2263), .ZN(n15605) );
NOR2_X1 U17680 ( .A1(n2271), .A2(n2272), .ZN(n2262) );
NOR2_X1 U17681 ( .A1(n2264), .A2(n2265), .ZN(n2263) );
NAND2_X1 U17682 ( .A1(n2273), .A2(n2274), .ZN(n2272) );
NAND2_X1 U17683 ( .A1(n2334), .A2(n2335), .ZN(n15593) );
NOR2_X1 U17684 ( .A1(n2358), .A2(n2359), .ZN(n2334) );
NOR2_X1 U17685 ( .A1(n2336), .A2(n2337), .ZN(n2335) );
NAND2_X1 U17686 ( .A1(n2360), .A2(n2361), .ZN(n2359) );
NAND2_X1 U17687 ( .A1(n2309), .A2(n2310), .ZN(n15604) );
NOR2_X1 U17688 ( .A1(n2320), .A2(n2321), .ZN(n2309) );
NOR2_X1 U17689 ( .A1(n2311), .A2(n2312), .ZN(n2310) );
NAND2_X1 U17690 ( .A1(n2109), .A2(n2322), .ZN(n2321) );
NAND2_X1 U17691 ( .A1(n2385), .A2(n2386), .ZN(n15574) );
AND2_X1 U17692 ( .A1(n2266), .A2(n2104), .ZN(n2386) );
NOR2_X1 U17693 ( .A1(n2389), .A2(n2390), .ZN(n2385) );
NOR2_X1 U17694 ( .A1(n16456), .A2(n2392), .ZN(n2389) );
NAND2_X1 U17695 ( .A1(n5185), .A2(n5186), .ZN(n15570) );
NOR2_X1 U17696 ( .A1(n5159), .A2(n5190), .ZN(n5185) );
NOR2_X1 U17697 ( .A1(n20987), .A2(n5188), .ZN(n5186) );
NAND2_X1 U17698 ( .A1(n5191), .A2(n5192), .ZN(n5190) );
INV_X1 U17699 ( .A(ex_block_i_alu_i_shift_amt_compl_0), .ZN(n20871) );
NOR2_X1 U17700 ( .A1(n5273), .A2(n20764), .ZN(n4257) );
INV_X1 U17701 ( .A(alu_operand_b_ex_2), .ZN(n20864) );
NAND2_X1 U17702 ( .A1(n9422), .A2(n9423), .ZN(n883) );
NOR2_X1 U17703 ( .A1(n9426), .A2(n9427), .ZN(n9422) );
NOR2_X1 U17704 ( .A1(n9424), .A2(n9425), .ZN(n9423) );
NOR2_X1 U17705 ( .A1(n8819), .A2(n15809), .ZN(n9426) );
NAND2_X1 U17706 ( .A1(n8865), .A2(n8866), .ZN(n323) );
NOR2_X1 U17707 ( .A1(n8869), .A2(n8870), .ZN(n8865) );
NOR2_X1 U17708 ( .A1(n8867), .A2(n8868), .ZN(n8866) );
NOR2_X1 U17709 ( .A1(n8819), .A2(n15806), .ZN(n8869) );
NAND2_X1 U17710 ( .A1(n8813), .A2(n8814), .ZN(n282) );
NOR2_X1 U17711 ( .A1(n8817), .A2(n8818), .ZN(n8813) );
NOR2_X1 U17712 ( .A1(n8815), .A2(n8816), .ZN(n8814) );
NOR2_X1 U17713 ( .A1(n8819), .A2(n15885), .ZN(n8817) );
INV_X1 U17714 ( .A(alu_operand_b_ex_1), .ZN(n20869) );
INV_X1 U17715 ( .A(alu_operand_b_ex_3), .ZN(n20861) );
NAND2_X1 U17716 ( .A1(n21023), .A2(n21022), .ZN(n21263) );
NAND2_X1 U17717 ( .A1(ex_block_i_alu_i_adder_in_a_2), .A2(n21229), .ZN(n21023) );
OR2_X1 U17718 ( .A1(n21229), .A2(ex_block_i_alu_i_adder_in_a_2), .ZN(n21021) );
NAND2_X1 U17719 ( .A1(n21032), .A2(n21031), .ZN(n21281) );
NAND2_X1 U17720 ( .A1(ex_block_i_alu_i_adder_in_a_5), .A2(n21275), .ZN(n21032) );
OR2_X1 U17721 ( .A1(n21275), .A2(ex_block_i_alu_i_adder_in_a_5), .ZN(n21030) );
NAND2_X1 U17722 ( .A1(n21035), .A2(n21034), .ZN(n21287) );
NAND2_X1 U17723 ( .A1(ex_block_i_alu_i_adder_in_a_6), .A2(n21281), .ZN(n21035) );
OR2_X1 U17724 ( .A1(n21281), .A2(ex_block_i_alu_i_adder_in_a_6), .ZN(n21033) );
NAND2_X1 U17725 ( .A1(n21044), .A2(n21043), .ZN(n21050) );
NAND2_X1 U17726 ( .A1(ex_block_i_alu_i_adder_in_a_9), .A2(n21299), .ZN(n21044) );
OR2_X1 U17727 ( .A1(n21299), .A2(ex_block_i_alu_i_adder_in_a_9), .ZN(n21042) );
NAND2_X1 U17728 ( .A1(n21053), .A2(n21052), .ZN(n21059) );
NAND2_X1 U17729 ( .A1(ex_block_i_alu_i_adder_in_a_10), .A2(n21050), .ZN(n21053) );
OR2_X1 U17730 ( .A1(n21050), .A2(ex_block_i_alu_i_adder_in_a_10), .ZN(n21051) );
NAND2_X1 U17731 ( .A1(n21071), .A2(n21070), .ZN(n21077) );
NAND2_X1 U17732 ( .A1(ex_block_i_alu_i_adder_in_a_12), .A2(n21068), .ZN(n21071) );
OR2_X1 U17733 ( .A1(n21068), .A2(ex_block_i_alu_i_adder_in_a_12), .ZN(n21069) );
INV_X1 U17734 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .ZN(n20789) );
INV_X1 U17735 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .ZN(n20792) );
INV_X1 U17736 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .ZN(n20786) );
INV_X1 U17737 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .ZN(n20795) );
INV_X1 U17738 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .ZN(n20783) );
INV_X1 U17739 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .ZN(n20798) );
INV_X1 U17740 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .ZN(n20780) );
INV_X1 U17741 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .ZN(n20801) );
INV_X1 U17742 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .ZN(n20777) );
INV_X1 U17743 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .ZN(n20774) );
INV_X1 U17744 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .ZN(n20771) );
INV_X1 U17745 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .ZN(n20768) );
INV_X1 U17746 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n20804) );
INV_X1 U17747 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n20765) );
INV_X1 U17748 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n20807) );
NOR2_X1 U17749 ( .A1(n8601), .A2(n20752), .ZN(n9887) );
NAND2_X1 U17750 ( .A1(n21020), .A2(n21019), .ZN(n21229) );
NAND2_X1 U17751 ( .A1(n20939), .A2(ex_block_i_alu_i_adder_in_a_1), .ZN(n21020) );
NAND2_X1 U17752 ( .A1(ex_block_i_alu_i_adder_in_b_1), .A2(n21018), .ZN(n21019) );
NAND2_X1 U17753 ( .A1(n16334), .A2(n20758), .ZN(n21018) );
NAND2_X1 U17754 ( .A1(n21029), .A2(n21028), .ZN(n21275) );
NAND2_X1 U17755 ( .A1(ex_block_i_alu_i_adder_in_a_4), .A2(n21269), .ZN(n21029) );
NAND2_X1 U17756 ( .A1(ex_block_i_alu_i_adder_in_b_4), .A2(n21027), .ZN(n21028) );
OR2_X1 U17757 ( .A1(n21269), .A2(ex_block_i_alu_i_adder_in_a_4), .ZN(n21027) );
NAND2_X1 U17758 ( .A1(n21038), .A2(n21037), .ZN(n21293) );
NAND2_X1 U17759 ( .A1(ex_block_i_alu_i_adder_in_a_7), .A2(n21287), .ZN(n21038) );
NAND2_X1 U17760 ( .A1(ex_block_i_alu_i_adder_in_b_7), .A2(n21036), .ZN(n21037) );
OR2_X1 U17761 ( .A1(n21287), .A2(ex_block_i_alu_i_adder_in_a_7), .ZN(n21036) );
NAND2_X1 U17762 ( .A1(n21041), .A2(n21040), .ZN(n21299) );
NAND2_X1 U17763 ( .A1(ex_block_i_alu_i_adder_in_a_8), .A2(n21293), .ZN(n21041) );
NAND2_X1 U17764 ( .A1(ex_block_i_alu_i_adder_in_b_8), .A2(n21039), .ZN(n21040) );
OR2_X1 U17765 ( .A1(n21293), .A2(ex_block_i_alu_i_adder_in_a_8), .ZN(n21039) );
NAND2_X1 U17766 ( .A1(n21062), .A2(n21061), .ZN(n21068) );
NAND2_X1 U17767 ( .A1(ex_block_i_alu_i_adder_in_a_11), .A2(n21059), .ZN(n21062) );
NAND2_X1 U17768 ( .A1(ex_block_i_alu_i_adder_in_b_11), .A2(n21060), .ZN(n21061) );
OR2_X1 U17769 ( .A1(n21059), .A2(ex_block_i_alu_i_adder_in_a_11), .ZN(n21060) );
NOR2_X1 U17770 ( .A1(n8601), .A2(n20756), .ZN(n9424) );
NOR2_X1 U17771 ( .A1(n16364), .A2(n20746), .ZN(n8867) );
NOR2_X1 U17772 ( .A1(n16364), .A2(n20741), .ZN(n8815) );
NAND2_X1 U17773 ( .A1(n6257), .A2(n6258), .ZN(ex_block_i_alu_i_adder_in_a_2) );
NAND2_X1 U17774 ( .A1(n6238), .A2(n15898), .ZN(n6257) );
NAND2_X1 U17775 ( .A1(n16357), .A2(n883), .ZN(n6258) );
NAND2_X1 U17776 ( .A1(n6245), .A2(n6246), .ZN(ex_block_i_alu_i_adder_in_a_5) );
NAND2_X1 U17777 ( .A1(n16408), .A2(n15901), .ZN(n6245) );
NAND2_X1 U17778 ( .A1(n16357), .A2(n282), .ZN(n6246) );
NAND2_X1 U17779 ( .A1(n6249), .A2(n6250), .ZN(ex_block_i_alu_i_adder_in_a_3) );
NAND2_X1 U17780 ( .A1(n16408), .A2(n15899), .ZN(n6249) );
NAND2_X1 U17781 ( .A1(n16357), .A2(n466), .ZN(n6250) );
NAND2_X1 U17782 ( .A1(n6247), .A2(n6248), .ZN(ex_block_i_alu_i_adder_in_a_4) );
NAND2_X1 U17783 ( .A1(n16408), .A2(n15900), .ZN(n6247) );
NAND2_X1 U17784 ( .A1(n20961), .A2(n323), .ZN(n6248) );
INV_X1 U17785 ( .A(n3437), .ZN(n19815) );
INV_X1 U17786 ( .A(n3432), .ZN(n19813) );
NAND2_X1 U17787 ( .A1(n21026), .A2(n21025), .ZN(n21269) );
NAND2_X1 U17788 ( .A1(ex_block_i_alu_i_adder_in_a_3), .A2(n21263), .ZN(n21026) );
OR2_X1 U17789 ( .A1(n21263), .A2(ex_block_i_alu_i_adder_in_a_3), .ZN(n21024) );
NAND2_X1 U17790 ( .A1(n6279), .A2(n6280), .ZN(ex_block_i_alu_i_adder_in_a_1) );
NAND2_X1 U17791 ( .A1(n6238), .A2(n15886), .ZN(n6280) );
NAND2_X1 U17792 ( .A1(n20961), .A2(n1391), .ZN(n6279) );
NOR2_X1 U17793 ( .A1(n394), .A2(n395), .ZN(n388) );
NOR2_X1 U17794 ( .A1(n83), .A2(n15857), .ZN(n395) );
NAND2_X1 U17795 ( .A1(n431), .A2(n432), .ZN(n423) );
NOR2_X1 U17796 ( .A1(n436), .A2(n437), .ZN(n431) );
NOR2_X1 U17797 ( .A1(n433), .A2(n434), .ZN(n432) );
NOR2_X1 U17798 ( .A1(n20818), .A2(n16208), .ZN(n437) );
NAND2_X1 U17799 ( .A1(n634), .A2(n635), .ZN(n626) );
NOR2_X1 U17800 ( .A1(n639), .A2(n640), .ZN(n634) );
NOR2_X1 U17801 ( .A1(n636), .A2(n637), .ZN(n635) );
NOR2_X1 U17802 ( .A1(n20818), .A2(n16241), .ZN(n640) );
NAND2_X1 U17803 ( .A1(n594), .A2(n595), .ZN(n586) );
NOR2_X1 U17804 ( .A1(n599), .A2(n600), .ZN(n594) );
NOR2_X1 U17805 ( .A1(n596), .A2(n597), .ZN(n595) );
NOR2_X1 U17806 ( .A1(n20818), .A2(n16244), .ZN(n600) );
NAND2_X1 U17807 ( .A1(n554), .A2(n555), .ZN(n546) );
NOR2_X1 U17808 ( .A1(n559), .A2(n560), .ZN(n554) );
NOR2_X1 U17809 ( .A1(n556), .A2(n557), .ZN(n555) );
NOR2_X1 U17810 ( .A1(n20818), .A2(n16202), .ZN(n560) );
NAND2_X1 U17811 ( .A1(n514), .A2(n515), .ZN(n506) );
NOR2_X1 U17812 ( .A1(n519), .A2(n520), .ZN(n514) );
NOR2_X1 U17813 ( .A1(n516), .A2(n517), .ZN(n515) );
NOR2_X1 U17814 ( .A1(n20818), .A2(n16205), .ZN(n520) );
NAND2_X1 U17815 ( .A1(n673), .A2(n674), .ZN(n665) );
NOR2_X1 U17816 ( .A1(n677), .A2(n678), .ZN(n673) );
NOR2_X1 U17817 ( .A1(n675), .A2(n676), .ZN(n674) );
NOR2_X1 U17818 ( .A1(n20818), .A2(n16238), .ZN(n678) );
NAND2_X1 U17819 ( .A1(n1343), .A2(n1344), .ZN(rf_wdata_wb_ecc_o_0_) );
NOR2_X1 U17820 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
NOR2_X1 U17821 ( .A1(n1376), .A2(n1377), .ZN(n1343) );
NAND2_X1 U17822 ( .A1(n1352), .A2(n1353), .ZN(n1345) );
NOR2_X1 U17823 ( .A1(n354), .A2(n355), .ZN(n353) );
NAND2_X1 U17824 ( .A1(n365), .A2(n366), .ZN(n354) );
NAND2_X1 U17825 ( .A1(n642), .A2(n643), .ZN(rf_wdata_wb_ecc_o_25_) );
NOR2_X1 U17826 ( .A1(n644), .A2(n645), .ZN(n643) );
NOR2_X1 U17827 ( .A1(n665), .A2(n666), .ZN(n642) );
NAND2_X1 U17828 ( .A1(n646), .A2(n647), .ZN(n645) );
NAND2_X1 U17829 ( .A1(n399), .A2(n400), .ZN(rf_wdata_wb_ecc_o_30_) );
NOR2_X1 U17830 ( .A1(n401), .A2(n402), .ZN(n400) );
NOR2_X1 U17831 ( .A1(n423), .A2(n424), .ZN(n399) );
NAND2_X1 U17832 ( .A1(n403), .A2(n404), .ZN(n402) );
NAND2_X1 U17833 ( .A1(n602), .A2(n603), .ZN(rf_wdata_wb_ecc_o_26_) );
NOR2_X1 U17834 ( .A1(n604), .A2(n605), .ZN(n603) );
NOR2_X1 U17835 ( .A1(n626), .A2(n627), .ZN(n602) );
NAND2_X1 U17836 ( .A1(n606), .A2(n607), .ZN(n605) );
NAND2_X1 U17837 ( .A1(n562), .A2(n563), .ZN(rf_wdata_wb_ecc_o_27_) );
NOR2_X1 U17838 ( .A1(n564), .A2(n565), .ZN(n563) );
NOR2_X1 U17839 ( .A1(n586), .A2(n587), .ZN(n562) );
NAND2_X1 U17840 ( .A1(n566), .A2(n567), .ZN(n565) );
NAND2_X1 U17841 ( .A1(n522), .A2(n523), .ZN(rf_wdata_wb_ecc_o_28_) );
NOR2_X1 U17842 ( .A1(n524), .A2(n525), .ZN(n523) );
NOR2_X1 U17843 ( .A1(n546), .A2(n547), .ZN(n522) );
NAND2_X1 U17844 ( .A1(n526), .A2(n527), .ZN(n525) );
NAND2_X1 U17845 ( .A1(n482), .A2(n483), .ZN(rf_wdata_wb_ecc_o_29_) );
NOR2_X1 U17846 ( .A1(n484), .A2(n485), .ZN(n483) );
NOR2_X1 U17847 ( .A1(n506), .A2(n507), .ZN(n482) );
NAND2_X1 U17848 ( .A1(n486), .A2(n487), .ZN(n485) );
INV_X1 U17849 ( .A(n197), .ZN(n20841) );
INV_X1 U17850 ( .A(n1297), .ZN(n20830) );
INV_X1 U17851 ( .A(n255), .ZN(n20846) );
NOR2_X1 U17852 ( .A1(n8601), .A2(n20711), .ZN(n9831) );
NOR2_X1 U17853 ( .A1(n16364), .A2(n20730), .ZN(n8728) );
NOR2_X1 U17854 ( .A1(n16364), .A2(n20724), .ZN(n8691) );
NOR2_X1 U17855 ( .A1(n16364), .A2(n20719), .ZN(n8639) );
NOR2_X1 U17856 ( .A1(n16364), .A2(n20715), .ZN(n8598) );
NOR2_X1 U17857 ( .A1(n16364), .A2(n20735), .ZN(n8771) );
NAND2_X1 U17858 ( .A1(n6243), .A2(n6244), .ZN(ex_block_i_alu_i_adder_in_a_6) );
NAND2_X1 U17859 ( .A1(n16408), .A2(n15902), .ZN(n6243) );
NAND2_X1 U17860 ( .A1(n16357), .A2(n240), .ZN(n6244) );
NAND2_X1 U17861 ( .A1(n6241), .A2(n6242), .ZN(ex_block_i_alu_i_adder_in_a_7) );
NAND2_X1 U17862 ( .A1(n16408), .A2(n15903), .ZN(n6241) );
NAND2_X1 U17863 ( .A1(n20961), .A2(n213), .ZN(n6242) );
NAND2_X1 U17864 ( .A1(n6239), .A2(n6240), .ZN(ex_block_i_alu_i_adder_in_a_8) );
NAND2_X1 U17865 ( .A1(n16408), .A2(n15904), .ZN(n6239) );
NAND2_X1 U17866 ( .A1(n16357), .A2(n170), .ZN(n6240) );
NAND2_X1 U17867 ( .A1(n6236), .A2(n6237), .ZN(ex_block_i_alu_i_adder_in_a_9) );
NAND2_X1 U17868 ( .A1(n16408), .A2(n15905), .ZN(n6236) );
NAND2_X1 U17869 ( .A1(n20961), .A2(n107), .ZN(n6237) );
NAND2_X1 U17870 ( .A1(n6297), .A2(n6298), .ZN(ex_block_i_alu_i_adder_in_a_11) );
NAND2_X1 U17871 ( .A1(n16408), .A2(n15896), .ZN(n6297) );
NAND2_X1 U17872 ( .A1(n20961), .A2(n1295), .ZN(n6298) );
INV_X1 U17873 ( .A(n3472), .ZN(n19831) );
INV_X1 U17874 ( .A(n3462), .ZN(n19826) );
INV_X1 U17875 ( .A(n3447), .ZN(n19818) );
NAND2_X1 U17876 ( .A1(n6299), .A2(n6300), .ZN(ex_block_i_alu_i_adder_in_a_10) );
NAND2_X1 U17877 ( .A1(n6238), .A2(n15906), .ZN(n6300) );
NAND2_X1 U17878 ( .A1(n16357), .A2(n51), .ZN(n6299) );
INV_X1 U17879 ( .A(n54), .ZN(n20833) );
INV_X1 U17880 ( .A(n109), .ZN(n20835) );
NAND2_X1 U17881 ( .A1(n3806), .A2(n3807), .ZN(n3467) );
NOR2_X1 U17882 ( .A1(n3777), .A2(n3813), .ZN(n3806) );
NOR2_X1 U17883 ( .A1(n3808), .A2(n3809), .ZN(n3807) );
NAND2_X1 U17884 ( .A1(n3814), .A2(n3815), .ZN(n3813) );
NAND2_X1 U17885 ( .A1(n3783), .A2(n3784), .ZN(n3457) );
NOR2_X1 U17886 ( .A1(n3777), .A2(n3790), .ZN(n3783) );
NOR2_X1 U17887 ( .A1(n3785), .A2(n3786), .ZN(n3784) );
NAND2_X1 U17888 ( .A1(n3791), .A2(n3792), .ZN(n3790) );
NAND2_X1 U17889 ( .A1(n3767), .A2(n3768), .ZN(n3452) );
NOR2_X1 U17890 ( .A1(n3777), .A2(n3778), .ZN(n3767) );
NOR2_X1 U17891 ( .A1(n3769), .A2(n3770), .ZN(n3768) );
NAND2_X1 U17892 ( .A1(n3779), .A2(n3780), .ZN(n3778) );
INV_X1 U17893 ( .A(n149), .ZN(n20839) );
NAND2_X1 U17894 ( .A1(n3810), .A2(n3811), .ZN(n3809) );
NAND2_X1 U17895 ( .A1(n3774), .A2(crash_dump_o_25_), .ZN(n3810) );
NAND2_X1 U17896 ( .A1(n3773), .A2(data_addr_o_25_), .ZN(n3811) );
NAND2_X1 U17897 ( .A1(n3787), .A2(n3788), .ZN(n3786) );
NAND2_X1 U17898 ( .A1(n3774), .A2(crash_dump_o_27_), .ZN(n3787) );
NAND2_X1 U17899 ( .A1(n3773), .A2(data_addr_o_27_), .ZN(n3788) );
NAND2_X1 U17900 ( .A1(n3771), .A2(n3772), .ZN(n3770) );
NAND2_X1 U17901 ( .A1(n3774), .A2(crash_dump_o_28_), .ZN(n3771) );
NAND2_X1 U17902 ( .A1(n3773), .A2(data_addr_o_28_), .ZN(n3772) );
NAND2_X1 U17903 ( .A1(n944), .A2(n945), .ZN(n936) );
NOR2_X1 U17904 ( .A1(n948), .A2(n949), .ZN(n944) );
NOR2_X1 U17905 ( .A1(n946), .A2(n947), .ZN(n945) );
NOR2_X1 U17906 ( .A1(n20818), .A2(n16211), .ZN(n949) );
NAND2_X1 U17907 ( .A1(n863), .A2(n864), .ZN(n855) );
NOR2_X1 U17908 ( .A1(n867), .A2(n868), .ZN(n863) );
NOR2_X1 U17909 ( .A1(n865), .A2(n866), .ZN(n864) );
NOR2_X1 U17910 ( .A1(n20818), .A2(n16214), .ZN(n868) );
NAND2_X1 U17911 ( .A1(n824), .A2(n825), .ZN(n816) );
NOR2_X1 U17912 ( .A1(n828), .A2(n829), .ZN(n824) );
NOR2_X1 U17913 ( .A1(n826), .A2(n827), .ZN(n825) );
NOR2_X1 U17914 ( .A1(n20818), .A2(n16232), .ZN(n829) );
NAND2_X1 U17915 ( .A1(n786), .A2(n787), .ZN(n778) );
NOR2_X1 U17916 ( .A1(n790), .A2(n791), .ZN(n786) );
NOR2_X1 U17917 ( .A1(n788), .A2(n789), .ZN(n787) );
NOR2_X1 U17918 ( .A1(n20818), .A2(n16235), .ZN(n791) );
NAND2_X1 U17919 ( .A1(n748), .A2(n749), .ZN(n740) );
NOR2_X1 U17920 ( .A1(n752), .A2(n753), .ZN(n748) );
NOR2_X1 U17921 ( .A1(n750), .A2(n751), .ZN(n749) );
NOR2_X1 U17922 ( .A1(n20818), .A2(n16217), .ZN(n753) );
NAND2_X1 U17923 ( .A1(n711), .A2(n712), .ZN(n703) );
NOR2_X1 U17924 ( .A1(n715), .A2(n716), .ZN(n711) );
NOR2_X1 U17925 ( .A1(n713), .A2(n714), .ZN(n712) );
NOR2_X1 U17926 ( .A1(n20818), .A2(n16220), .ZN(n716) );
NAND2_X1 U17927 ( .A1(n913), .A2(n914), .ZN(rf_wdata_wb_ecc_o_19_) );
NOR2_X1 U17928 ( .A1(n915), .A2(n916), .ZN(n914) );
NOR2_X1 U17929 ( .A1(n936), .A2(n937), .ZN(n913) );
NAND2_X1 U17930 ( .A1(n917), .A2(n918), .ZN(n916) );
NAND2_X1 U17931 ( .A1(n832), .A2(n833), .ZN(rf_wdata_wb_ecc_o_20_) );
NOR2_X1 U17932 ( .A1(n834), .A2(n835), .ZN(n833) );
NOR2_X1 U17933 ( .A1(n855), .A2(n856), .ZN(n832) );
NAND2_X1 U17934 ( .A1(n836), .A2(n837), .ZN(n835) );
NAND2_X1 U17935 ( .A1(n793), .A2(n794), .ZN(rf_wdata_wb_ecc_o_21_) );
NOR2_X1 U17936 ( .A1(n795), .A2(n796), .ZN(n794) );
NOR2_X1 U17937 ( .A1(n816), .A2(n817), .ZN(n793) );
NAND2_X1 U17938 ( .A1(n797), .A2(n798), .ZN(n796) );
NAND2_X1 U17939 ( .A1(n755), .A2(n756), .ZN(rf_wdata_wb_ecc_o_22_) );
NOR2_X1 U17940 ( .A1(n757), .A2(n758), .ZN(n756) );
NOR2_X1 U17941 ( .A1(n778), .A2(n779), .ZN(n755) );
NAND2_X1 U17942 ( .A1(n759), .A2(n760), .ZN(n758) );
NAND2_X1 U17943 ( .A1(n718), .A2(n719), .ZN(rf_wdata_wb_ecc_o_23_) );
NOR2_X1 U17944 ( .A1(n720), .A2(n721), .ZN(n719) );
NOR2_X1 U17945 ( .A1(n740), .A2(n741), .ZN(n718) );
NAND2_X1 U17946 ( .A1(n722), .A2(n723), .ZN(n721) );
NAND2_X1 U17947 ( .A1(n680), .A2(n681), .ZN(rf_wdata_wb_ecc_o_24_) );
NOR2_X1 U17948 ( .A1(n682), .A2(n683), .ZN(n681) );
NOR2_X1 U17949 ( .A1(n703), .A2(n704), .ZN(n680) );
NAND2_X1 U17950 ( .A1(n684), .A2(n685), .ZN(n683) );
NAND2_X1 U17951 ( .A1(n6146), .A2(n6147), .ZN(n6145) );
NAND2_X1 U17952 ( .A1(n16410), .A2(n20691), .ZN(n6147) );
NAND2_X1 U17953 ( .A1(n5916), .A2(n20811), .ZN(n6146) );
NOR2_X1 U17954 ( .A1(n359), .A2(n20207), .ZN(n516) );
NOR2_X1 U17955 ( .A1(n359), .A2(n20169), .ZN(n433) );
NOR2_X1 U17956 ( .A1(n92), .A2(n20207), .ZN(n1202) );
NOR2_X1 U17957 ( .A1(n92), .A2(n20169), .ZN(n1163) );
NOR2_X1 U17958 ( .A1(n92), .A2(n20107), .ZN(n1124) );
NOR2_X1 U17959 ( .A1(n8601), .A2(n20695), .ZN(n9669) );
NOR2_X1 U17960 ( .A1(n16364), .A2(n20699), .ZN(n9706) );
NOR2_X1 U17961 ( .A1(n8601), .A2(n20703), .ZN(n9746) );
NOR2_X1 U17962 ( .A1(n16364), .A2(n20707), .ZN(n9794) );
NOR2_X1 U17963 ( .A1(n8601), .A2(n20687), .ZN(n9594) );
NOR2_X1 U17964 ( .A1(n8601), .A2(n20691), .ZN(n9632) );
NAND2_X1 U17965 ( .A1(n6122), .A2(n6123), .ZN(ex_block_i_alu_i_adder_in_b_17) );
NOR2_X1 U17966 ( .A1(n6131), .A2(n6132), .ZN(n6122) );
NOR2_X1 U17967 ( .A1(n6124), .A2(n6125), .ZN(n6123) );
NOR2_X1 U17968 ( .A1(n5917), .A2(n16109), .ZN(n6131) );
NAND2_X1 U17969 ( .A1(n6295), .A2(n6296), .ZN(ex_block_i_alu_i_adder_in_a_12) );
NAND2_X1 U17970 ( .A1(n16408), .A2(n15897), .ZN(n6295) );
NAND2_X1 U17971 ( .A1(n20961), .A2(n1258), .ZN(n6296) );
NAND2_X1 U17972 ( .A1(n6293), .A2(n6294), .ZN(ex_block_i_alu_i_adder_in_a_13) );
NAND2_X1 U17973 ( .A1(n6238), .A2(n15880), .ZN(n6293) );
NAND2_X1 U17974 ( .A1(n20961), .A2(n1217), .ZN(n6294) );
NAND2_X1 U17975 ( .A1(n6291), .A2(n6292), .ZN(ex_block_i_alu_i_adder_in_a_14) );
NAND2_X1 U17976 ( .A1(n16408), .A2(n15881), .ZN(n6291) );
NAND2_X1 U17977 ( .A1(n20961), .A2(n1178), .ZN(n6292) );
NAND2_X1 U17978 ( .A1(n6289), .A2(n6290), .ZN(ex_block_i_alu_i_adder_in_a_15) );
NAND2_X1 U17979 ( .A1(n6238), .A2(n15882), .ZN(n6289) );
NAND2_X1 U17980 ( .A1(n20961), .A2(n1139), .ZN(n6290) );
NAND2_X1 U17981 ( .A1(n6287), .A2(n6288), .ZN(ex_block_i_alu_i_adder_in_a_16) );
NAND2_X1 U17982 ( .A1(n16408), .A2(n15883), .ZN(n6287) );
NAND2_X1 U17983 ( .A1(n20961), .A2(n1102), .ZN(n6288) );
NAND2_X1 U17984 ( .A1(n6285), .A2(n6286), .ZN(ex_block_i_alu_i_adder_in_a_17) );
NAND2_X1 U17985 ( .A1(n6238), .A2(n15861), .ZN(n6285) );
NAND2_X1 U17986 ( .A1(n20961), .A2(n1046), .ZN(n6286) );
INV_X1 U17987 ( .A(n3513), .ZN(n19846) );
INV_X1 U17988 ( .A(n3508), .ZN(n19843) );
INV_X1 U17989 ( .A(n3487), .ZN(n19838) );
INV_X1 U17990 ( .A(n3482), .ZN(n19836) );
INV_X1 U17991 ( .A(n3477), .ZN(n19833) );
NAND2_X1 U17992 ( .A1(n1029), .A2(n1030), .ZN(rf_wdata_wb_ecc_o_16_) );
NOR2_X1 U17993 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U17994 ( .A1(n1071), .A2(n1072), .ZN(n1029) );
NAND2_X1 U17995 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U17996 ( .A1(n6162), .A2(n6163), .ZN(ex_block_i_alu_i_adder_in_b_14) );
NOR2_X1 U17997 ( .A1(n6172), .A2(n6173), .ZN(n6162) );
NOR2_X1 U17998 ( .A1(n6164), .A2(n6165), .ZN(n6163) );
NOR2_X1 U17999 ( .A1(n5917), .A2(n16112), .ZN(n6172) );
INV_X1 U18000 ( .A(n1256), .ZN(n20828) );
NAND2_X1 U18001 ( .A1(n6193), .A2(n6194), .ZN(n6192) );
NAND2_X1 U18002 ( .A1(n16410), .A2(n20703), .ZN(n6194) );
NAND2_X1 U18003 ( .A1(n5916), .A2(n20817), .ZN(n6193) );
NAND2_X1 U18004 ( .A1(n6174), .A2(n6175), .ZN(n6173) );
NAND2_X1 U18005 ( .A1(n16410), .A2(n20699), .ZN(n6175) );
NAND2_X1 U18006 ( .A1(n5916), .A2(n20815), .ZN(n6174) );
NAND2_X1 U18007 ( .A1(n6160), .A2(n6161), .ZN(n6159) );
NAND2_X1 U18008 ( .A1(n16410), .A2(n20695), .ZN(n6161) );
NAND2_X1 U18009 ( .A1(n5916), .A2(n20813), .ZN(n6160) );
NAND2_X1 U18010 ( .A1(n3862), .A2(n3863), .ZN(n3492) );
NOR2_X1 U18011 ( .A1(n3777), .A2(n3869), .ZN(n3862) );
NOR2_X1 U18012 ( .A1(n3864), .A2(n3865), .ZN(n3863) );
NAND2_X1 U18013 ( .A1(n3870), .A2(n3871), .ZN(n3869) );
NAND2_X1 U18014 ( .A1(n6176), .A2(n6177), .ZN(ex_block_i_alu_i_adder_in_b_13) );
NOR2_X1 U18015 ( .A1(n6191), .A2(n6192), .ZN(n6176) );
NOR2_X1 U18016 ( .A1(n6178), .A2(n6179), .ZN(n6177) );
NOR2_X1 U18017 ( .A1(n5917), .A2(n16113), .ZN(n6191) );
NAND2_X1 U18018 ( .A1(n6148), .A2(n6149), .ZN(ex_block_i_alu_i_adder_in_b_15) );
NOR2_X1 U18019 ( .A1(n6158), .A2(n6159), .ZN(n6148) );
NOR2_X1 U18020 ( .A1(n6150), .A2(n6151), .ZN(n6149) );
NOR2_X1 U18021 ( .A1(n5917), .A2(n16111), .ZN(n6158) );
NAND2_X1 U18022 ( .A1(n6135), .A2(n6136), .ZN(ex_block_i_alu_i_adder_in_b_16) );
NOR2_X1 U18023 ( .A1(n6144), .A2(n6145), .ZN(n6135) );
NOR2_X1 U18024 ( .A1(n6137), .A2(n6138), .ZN(n6136) );
NOR2_X1 U18025 ( .A1(n5917), .A2(n16110), .ZN(n6144) );
NAND2_X1 U18026 ( .A1(n6139), .A2(n6140), .ZN(n6138) );
NAND2_X1 U18027 ( .A1(n1100), .A2(n5904), .ZN(n6139) );
NAND2_X1 U18028 ( .A1(n20810), .A2(n5826), .ZN(n6140) );
NAND2_X1 U18029 ( .A1(n6126), .A2(n6127), .ZN(n6125) );
NAND2_X1 U18030 ( .A1(n1044), .A2(n5904), .ZN(n6126) );
NAND2_X1 U18031 ( .A1(n20808), .A2(n5826), .ZN(n6127) );
INV_X1 U18032 ( .A(n1100), .ZN(n20810) );
INV_X1 U18033 ( .A(n1044), .ZN(n20808) );
NAND2_X1 U18034 ( .A1(n3866), .A2(n3867), .ZN(n3865) );
NAND2_X1 U18035 ( .A1(n3774), .A2(crash_dump_o_20_), .ZN(n3866) );
NAND2_X1 U18036 ( .A1(n3773), .A2(data_addr_o_20_), .ZN(n3867) );
NAND2_X1 U18037 ( .A1(n6180), .A2(n6181), .ZN(n6179) );
NAND2_X1 U18038 ( .A1(n1219), .A2(n5904), .ZN(n6180) );
NAND2_X1 U18039 ( .A1(n20816), .A2(n16409), .ZN(n6181) );
INV_X1 U18040 ( .A(n1219), .ZN(n20816) );
NAND2_X1 U18041 ( .A1(n6166), .A2(n6167), .ZN(n6165) );
NAND2_X1 U18042 ( .A1(n1180), .A2(n16334), .ZN(n6166) );
NAND2_X1 U18043 ( .A1(n20814), .A2(n5826), .ZN(n6167) );
INV_X1 U18044 ( .A(n1180), .ZN(n20814) );
NAND2_X1 U18045 ( .A1(n6152), .A2(n6153), .ZN(n6151) );
NAND2_X1 U18046 ( .A1(n1141), .A2(n5904), .ZN(n6152) );
NAND2_X1 U18047 ( .A1(n20812), .A2(n5826), .ZN(n6153) );
INV_X1 U18048 ( .A(n1141), .ZN(n20812) );
NAND2_X1 U18049 ( .A1(n356), .A2(n357), .ZN(n355) );
NOR2_X1 U18050 ( .A1(n360), .A2(n361), .ZN(n356) );
OR2_X1 U18051 ( .A1(n20107), .A2(n359), .ZN(n357) );
NOR2_X1 U18052 ( .A1(n20014), .A2(n363), .ZN(n361) );
NAND2_X1 U18053 ( .A1(n1079), .A2(n1080), .ZN(n1071) );
NOR2_X1 U18054 ( .A1(n1084), .A2(n1085), .ZN(n1079) );
NOR2_X1 U18055 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U18056 ( .A1(n20818), .A2(n16223), .ZN(n1085) );
NAND2_X1 U18057 ( .A1(n1021), .A2(n1022), .ZN(n1013) );
NOR2_X1 U18058 ( .A1(n1025), .A2(n1026), .ZN(n1021) );
NOR2_X1 U18059 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NOR2_X1 U18060 ( .A1(n20818), .A2(n16226), .ZN(n1026) );
NAND2_X1 U18061 ( .A1(n983), .A2(n984), .ZN(n975) );
NOR2_X1 U18062 ( .A1(n987), .A2(n988), .ZN(n983) );
NOR2_X1 U18063 ( .A1(n985), .A2(n986), .ZN(n984) );
NOR2_X1 U18064 ( .A1(n20818), .A2(n16229), .ZN(n988) );
NAND2_X1 U18065 ( .A1(n1127), .A2(n1128), .ZN(rf_wdata_wb_ecc_o_14_) );
NOR2_X1 U18066 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U18067 ( .A1(n1154), .A2(n1155), .ZN(n1127) );
NAND2_X1 U18068 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U18069 ( .A1(n991), .A2(n992), .ZN(rf_wdata_wb_ecc_o_17_) );
NOR2_X1 U18070 ( .A1(n993), .A2(n994), .ZN(n992) );
NOR2_X1 U18071 ( .A1(n1013), .A2(n1014), .ZN(n991) );
NAND2_X1 U18072 ( .A1(n995), .A2(n996), .ZN(n994) );
NAND2_X1 U18073 ( .A1(n952), .A2(n953), .ZN(rf_wdata_wb_ecc_o_18_) );
NOR2_X1 U18074 ( .A1(n954), .A2(n955), .ZN(n953) );
NOR2_X1 U18075 ( .A1(n975), .A2(n976), .ZN(n952) );
NAND2_X1 U18076 ( .A1(n956), .A2(n957), .ZN(n955) );
NAND2_X1 U18077 ( .A1(n1166), .A2(n1167), .ZN(rf_wdata_wb_ecc_o_13_) );
NOR2_X1 U18078 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NOR2_X1 U18079 ( .A1(n1193), .A2(n1194), .ZN(n1166) );
NAND2_X1 U18080 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NAND2_X1 U18081 ( .A1(n1088), .A2(n1089), .ZN(rf_wdata_wb_ecc_o_15_) );
NOR2_X1 U18082 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U18083 ( .A1(n1115), .A2(n1116), .ZN(n1088) );
NAND2_X1 U18084 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U18085 ( .A1(n6133), .A2(n6134), .ZN(n6132) );
NAND2_X1 U18086 ( .A1(n16410), .A2(n20687), .ZN(n6134) );
NAND2_X1 U18087 ( .A1(n5916), .A2(n20809), .ZN(n6133) );
NAND2_X1 U18088 ( .A1(n6120), .A2(n6121), .ZN(n6119) );
NAND2_X1 U18089 ( .A1(n16410), .A2(n20680), .ZN(n6121) );
NAND2_X1 U18090 ( .A1(n5916), .A2(n20806), .ZN(n6120) );
NAND2_X1 U18091 ( .A1(n6106), .A2(n6107), .ZN(n6105) );
NAND2_X1 U18092 ( .A1(n16410), .A2(n20646), .ZN(n6107) );
NAND2_X1 U18093 ( .A1(n5916), .A2(n20803), .ZN(n6106) );
NAND2_X1 U18094 ( .A1(n6082), .A2(n6083), .ZN(n6081) );
NAND2_X1 U18095 ( .A1(n16410), .A2(n20608), .ZN(n6083) );
NAND2_X1 U18096 ( .A1(n5916), .A2(n20800), .ZN(n6082) );
NAND2_X1 U18097 ( .A1(n6066), .A2(n6067), .ZN(n6065) );
NAND2_X1 U18098 ( .A1(n5818), .A2(n20568), .ZN(n6067) );
NAND2_X1 U18099 ( .A1(n5916), .A2(n20797), .ZN(n6066) );
NAND2_X1 U18100 ( .A1(n6052), .A2(n6053), .ZN(n6051) );
NAND2_X1 U18101 ( .A1(n5818), .A2(n20528), .ZN(n6053) );
NAND2_X1 U18102 ( .A1(n5916), .A2(n20794), .ZN(n6052) );
NOR2_X1 U18103 ( .A1(n359), .A2(n20320), .ZN(n636) );
NOR2_X1 U18104 ( .A1(n359), .A2(n20283), .ZN(n596) );
NOR2_X1 U18105 ( .A1(n359), .A2(n20245), .ZN(n556) );
NOR2_X1 U18106 ( .A1(n92), .A2(n20357), .ZN(n88) );
NOR2_X1 U18107 ( .A1(n92), .A2(n20320), .ZN(n1339) );
NOR2_X1 U18108 ( .A1(n92), .A2(n20283), .ZN(n1280) );
NOR2_X1 U18109 ( .A1(n92), .A2(n20245), .ZN(n1241) );
NOR2_X1 U18110 ( .A1(n20357), .A2(n359), .ZN(n675) );
INV_X1 U18111 ( .A(n5104), .ZN(n20085) );
NOR2_X1 U18112 ( .A1(n8601), .A2(n20488), .ZN(n9296) );
NOR2_X1 U18113 ( .A1(n8601), .A2(n20568), .ZN(n9381) );
NOR2_X1 U18114 ( .A1(n8601), .A2(n20608), .ZN(n9467) );
NOR2_X1 U18115 ( .A1(n8601), .A2(n20646), .ZN(n9508) );
NOR2_X1 U18116 ( .A1(n8601), .A2(n20528), .ZN(n9339) );
NOR2_X1 U18117 ( .A1(n8601), .A2(n20680), .ZN(n9552) );
NAND2_X1 U18118 ( .A1(n6108), .A2(n6109), .ZN(ex_block_i_alu_i_adder_in_b_18) );
NOR2_X1 U18119 ( .A1(n6118), .A2(n6119), .ZN(n6108) );
NOR2_X1 U18120 ( .A1(n6110), .A2(n6111), .ZN(n6109) );
NOR2_X1 U18121 ( .A1(n5917), .A2(n16108), .ZN(n6118) );
NAND2_X1 U18122 ( .A1(n6054), .A2(n6055), .ZN(ex_block_i_alu_i_adder_in_b_21) );
NOR2_X1 U18123 ( .A1(n6064), .A2(n6065), .ZN(n6054) );
NOR2_X1 U18124 ( .A1(n6056), .A2(n6057), .ZN(n6055) );
NOR2_X1 U18125 ( .A1(n5917), .A2(n16105), .ZN(n6064) );
NAND2_X1 U18126 ( .A1(n6277), .A2(n6278), .ZN(ex_block_i_alu_i_adder_in_a_20) );
NAND2_X1 U18127 ( .A1(n16408), .A2(n15864), .ZN(n6277) );
NAND2_X1 U18128 ( .A1(n16357), .A2(n926), .ZN(n6278) );
NAND2_X1 U18129 ( .A1(n6275), .A2(n6276), .ZN(ex_block_i_alu_i_adder_in_a_21) );
NAND2_X1 U18130 ( .A1(n6238), .A2(n15865), .ZN(n6275) );
NAND2_X1 U18131 ( .A1(n16357), .A2(n845), .ZN(n6276) );
NAND2_X1 U18132 ( .A1(n6271), .A2(n6272), .ZN(ex_block_i_alu_i_adder_in_a_23) );
NAND2_X1 U18133 ( .A1(n6238), .A2(n15867), .ZN(n6271) );
NAND2_X1 U18134 ( .A1(n16357), .A2(n768), .ZN(n6272) );
NAND2_X1 U18135 ( .A1(n6273), .A2(n6274), .ZN(ex_block_i_alu_i_adder_in_a_22) );
NAND2_X1 U18136 ( .A1(n6238), .A2(n15866), .ZN(n6273) );
NAND2_X1 U18137 ( .A1(n16357), .A2(n806), .ZN(n6274) );
INV_X1 U18138 ( .A(n3543), .ZN(n19861) );
INV_X1 U18139 ( .A(n3538), .ZN(n19858) );
INV_X1 U18140 ( .A(n3533), .ZN(n19856) );
INV_X1 U18141 ( .A(n3528), .ZN(n19853) );
INV_X1 U18142 ( .A(n3518), .ZN(n19848) );
NAND2_X1 U18143 ( .A1(n3907), .A2(n3908), .ZN(n3523) );
NOR2_X1 U18144 ( .A1(n3777), .A2(n3914), .ZN(n3907) );
NOR2_X1 U18145 ( .A1(n3909), .A2(n3910), .ZN(n3908) );
NAND2_X1 U18146 ( .A1(n3915), .A2(n3916), .ZN(n3914) );
NAND2_X1 U18147 ( .A1(n6283), .A2(n6284), .ZN(ex_block_i_alu_i_adder_in_a_18) );
NAND2_X1 U18148 ( .A1(n6238), .A2(n15862), .ZN(n6283) );
NAND2_X1 U18149 ( .A1(n20961), .A2(n1003), .ZN(n6284) );
NAND2_X1 U18150 ( .A1(n6281), .A2(n6282), .ZN(ex_block_i_alu_i_adder_in_a_19) );
NAND2_X1 U18151 ( .A1(n16408), .A2(n15863), .ZN(n6281) );
NAND2_X1 U18152 ( .A1(n20961), .A2(n965), .ZN(n6282) );
NAND2_X1 U18153 ( .A1(n6094), .A2(n6095), .ZN(ex_block_i_alu_i_adder_in_b_19) );
NOR2_X1 U18154 ( .A1(n6104), .A2(n6105), .ZN(n6094) );
NOR2_X1 U18155 ( .A1(n6096), .A2(n6097), .ZN(n6095) );
NOR2_X1 U18156 ( .A1(n5917), .A2(n16107), .ZN(n6104) );
NAND2_X1 U18157 ( .A1(n6068), .A2(n6069), .ZN(ex_block_i_alu_i_adder_in_b_20) );
NOR2_X1 U18158 ( .A1(n6080), .A2(n6081), .ZN(n6068) );
NOR2_X1 U18159 ( .A1(n6070), .A2(n6071), .ZN(n6069) );
NOR2_X1 U18160 ( .A1(n5917), .A2(n16106), .ZN(n6080) );
NAND2_X1 U18161 ( .A1(n6040), .A2(n6041), .ZN(ex_block_i_alu_i_adder_in_b_22) );
NOR2_X1 U18162 ( .A1(n6050), .A2(n6051), .ZN(n6040) );
NOR2_X1 U18163 ( .A1(n6042), .A2(n6043), .ZN(n6041) );
NOR2_X1 U18164 ( .A1(n5917), .A2(n16104), .ZN(n6050) );
NAND2_X1 U18165 ( .A1(n6026), .A2(n6027), .ZN(ex_block_i_alu_i_adder_in_b_23) );
NOR2_X1 U18166 ( .A1(n6036), .A2(n6037), .ZN(n6026) );
NOR2_X1 U18167 ( .A1(n6028), .A2(n6029), .ZN(n6027) );
NOR2_X1 U18168 ( .A1(n5917), .A2(n16103), .ZN(n6036) );
NAND2_X1 U18169 ( .A1(n6112), .A2(n6113), .ZN(n6111) );
NAND2_X1 U18170 ( .A1(n1005), .A2(n16334), .ZN(n6112) );
NAND2_X1 U18171 ( .A1(n20805), .A2(n5826), .ZN(n6113) );
INV_X1 U18172 ( .A(n1005), .ZN(n20805) );
NAND2_X1 U18173 ( .A1(n6098), .A2(n6099), .ZN(n6097) );
NAND2_X1 U18174 ( .A1(n967), .A2(n16334), .ZN(n6098) );
NAND2_X1 U18175 ( .A1(n20802), .A2(n5826), .ZN(n6099) );
INV_X1 U18176 ( .A(n967), .ZN(n20802) );
NAND2_X1 U18177 ( .A1(n6072), .A2(n6073), .ZN(n6071) );
NAND2_X1 U18178 ( .A1(n928), .A2(n16334), .ZN(n6072) );
NAND2_X1 U18179 ( .A1(n20799), .A2(n16409), .ZN(n6073) );
INV_X1 U18180 ( .A(n928), .ZN(n20799) );
NAND2_X1 U18181 ( .A1(n6058), .A2(n6059), .ZN(n6057) );
NAND2_X1 U18182 ( .A1(n847), .A2(n16334), .ZN(n6058) );
NAND2_X1 U18183 ( .A1(n20796), .A2(n5826), .ZN(n6059) );
INV_X1 U18184 ( .A(n847), .ZN(n20796) );
NAND2_X1 U18185 ( .A1(n6044), .A2(n6045), .ZN(n6043) );
NAND2_X1 U18186 ( .A1(n808), .A2(n5904), .ZN(n6044) );
NAND2_X1 U18187 ( .A1(n20793), .A2(n16409), .ZN(n6045) );
INV_X1 U18188 ( .A(n808), .ZN(n20793) );
NAND2_X1 U18189 ( .A1(n6030), .A2(n6031), .ZN(n6029) );
NAND2_X1 U18190 ( .A1(n770), .A2(n5904), .ZN(n6030) );
NAND2_X1 U18191 ( .A1(n20790), .A2(n5826), .ZN(n6031) );
INV_X1 U18192 ( .A(n770), .ZN(n20790) );
NAND2_X1 U18193 ( .A1(n3911), .A2(n3912), .ZN(n3910) );
NAND2_X1 U18194 ( .A1(n3774), .A2(crash_dump_o_16_), .ZN(n3911) );
NAND2_X1 U18195 ( .A1(n3773), .A2(data_addr_o_16_), .ZN(n3912) );
NAND2_X1 U18196 ( .A1(n34), .A2(n35), .ZN(rf_wdata_wb_ecc_o_9_) );
NOR2_X1 U18197 ( .A1(n36), .A2(n37), .ZN(n35) );
NOR2_X1 U18198 ( .A1(n74), .A2(n75), .ZN(n34) );
NAND2_X1 U18199 ( .A1(n38), .A2(n39), .ZN(n37) );
NAND2_X1 U18200 ( .A1(n1283), .A2(n1284), .ZN(rf_wdata_wb_ecc_o_10_) );
NOR2_X1 U18201 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NOR2_X1 U18202 ( .A1(n1327), .A2(n1328), .ZN(n1283) );
NAND2_X1 U18203 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
NAND2_X1 U18204 ( .A1(n1244), .A2(n1245), .ZN(rf_wdata_wb_ecc_o_11_) );
NOR2_X1 U18205 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
NOR2_X1 U18206 ( .A1(n1271), .A2(n1272), .ZN(n1244) );
NAND2_X1 U18207 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND2_X1 U18208 ( .A1(n1205), .A2(n1206), .ZN(rf_wdata_wb_ecc_o_12_) );
NOR2_X1 U18209 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NOR2_X1 U18210 ( .A1(n1232), .A2(n1233), .ZN(n1205) );
NAND2_X1 U18211 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NOR2_X1 U18212 ( .A1(n20869), .A2(ex_block_i_alu_i_shift_amt_compl_0), .ZN(n7719) );
NAND2_X1 U18213 ( .A1(n6038), .A2(n6039), .ZN(n6037) );
NAND2_X1 U18214 ( .A1(n5818), .A2(n20488), .ZN(n6039) );
NAND2_X1 U18215 ( .A1(n5916), .A2(n20791), .ZN(n6038) );
NAND2_X1 U18216 ( .A1(n6024), .A2(n6025), .ZN(n6023) );
NAND2_X1 U18217 ( .A1(n5818), .A2(n20448), .ZN(n6025) );
NAND2_X1 U18218 ( .A1(n5916), .A2(n20788), .ZN(n6024) );
NAND2_X1 U18219 ( .A1(n6010), .A2(n6011), .ZN(n6009) );
NAND2_X1 U18220 ( .A1(n16410), .A2(n20408), .ZN(n6011) );
NAND2_X1 U18221 ( .A1(n5916), .A2(n20785), .ZN(n6010) );
NAND2_X1 U18222 ( .A1(n5996), .A2(n5997), .ZN(n5995) );
NAND2_X1 U18223 ( .A1(n5818), .A2(n20369), .ZN(n5997) );
NAND2_X1 U18224 ( .A1(n5916), .A2(n20782), .ZN(n5996) );
NAND2_X1 U18225 ( .A1(n5982), .A2(n5983), .ZN(n5981) );
NAND2_X1 U18226 ( .A1(n16410), .A2(n20330), .ZN(n5983) );
NAND2_X1 U18227 ( .A1(n5916), .A2(n20779), .ZN(n5982) );
NAND2_X1 U18228 ( .A1(n5968), .A2(n5969), .ZN(n5967) );
NAND2_X1 U18229 ( .A1(n5818), .A2(n20291), .ZN(n5969) );
NAND2_X1 U18230 ( .A1(n5916), .A2(n20776), .ZN(n5968) );
NOR2_X1 U18231 ( .A1(n10001), .A2(n9841), .ZN(n8106) );
NAND2_X1 U18232 ( .A1(n1297), .A2(n10002), .ZN(n10001) );
NAND2_X1 U18233 ( .A1(n1432), .A2(n149), .ZN(n9970) );
NAND2_X1 U18234 ( .A1(n1432), .A2(n1256), .ZN(n10002) );
NOR2_X1 U18235 ( .A1(n92), .A2(n20507), .ZN(n266) );
NOR2_X1 U18236 ( .A1(n92), .A2(n20469), .ZN(n224) );
NOR2_X1 U18237 ( .A1(n92), .A2(n20431), .ZN(n181) );
NOR2_X1 U18238 ( .A1(n92), .A2(n20394), .ZN(n133) );
NAND2_X1 U18239 ( .A1(n10346), .A2(n7678), .ZN(n7657) );
AND2_X1 U18240 ( .A1(n7623), .A2(n7622), .ZN(n10346) );
NAND2_X1 U18241 ( .A1(n1432), .A2(n255), .ZN(n10043) );
NOR2_X1 U18242 ( .A1(n20507), .A2(n359), .ZN(n826) );
NOR2_X1 U18243 ( .A1(n20469), .A2(n359), .ZN(n788) );
NOR2_X1 U18244 ( .A1(n20431), .A2(n359), .ZN(n750) );
NOR2_X1 U18245 ( .A1(n20394), .A2(n359), .ZN(n713) );
INV_X1 U18246 ( .A(n8056), .ZN(n20880) );
NOR2_X1 U18247 ( .A1(n367), .A2(n368), .ZN(n366) );
NOR2_X1 U18248 ( .A1(n20761), .A2(n370), .ZN(n368) );
NOR2_X1 U18249 ( .A1(n371), .A2(n15795), .ZN(n370) );
NOR2_X1 U18250 ( .A1(n20136), .A2(n15794), .ZN(n371) );
NAND2_X1 U18251 ( .A1(n923), .A2(n924), .ZN(n915) );
NOR2_X1 U18252 ( .A1(n929), .A2(n930), .ZN(n923) );
NOR2_X1 U18253 ( .A1(n367), .A2(n925), .ZN(n924) );
NOR2_X1 U18254 ( .A1(n20010), .A2(n378), .ZN(n930) );
NAND2_X1 U18255 ( .A1(n842), .A2(n843), .ZN(n834) );
NOR2_X1 U18256 ( .A1(n848), .A2(n849), .ZN(n842) );
NOR2_X1 U18257 ( .A1(n367), .A2(n844), .ZN(n843) );
NOR2_X1 U18258 ( .A1(n20009), .A2(n378), .ZN(n849) );
NAND2_X1 U18259 ( .A1(n803), .A2(n804), .ZN(n795) );
NOR2_X1 U18260 ( .A1(n809), .A2(n810), .ZN(n803) );
NOR2_X1 U18261 ( .A1(n367), .A2(n805), .ZN(n804) );
NOR2_X1 U18262 ( .A1(n20008), .A2(n378), .ZN(n810) );
NAND2_X1 U18263 ( .A1(n765), .A2(n766), .ZN(n757) );
NOR2_X1 U18264 ( .A1(n771), .A2(n772), .ZN(n765) );
NOR2_X1 U18265 ( .A1(n367), .A2(n767), .ZN(n766) );
NOR2_X1 U18266 ( .A1(n20007), .A2(n378), .ZN(n772) );
NAND2_X1 U18267 ( .A1(n727), .A2(n728), .ZN(n720) );
NOR2_X1 U18268 ( .A1(n733), .A2(n734), .ZN(n727) );
NOR2_X1 U18269 ( .A1(n367), .A2(n729), .ZN(n728) );
NOR2_X1 U18270 ( .A1(n20006), .A2(n378), .ZN(n734) );
NAND2_X1 U18271 ( .A1(n690), .A2(n691), .ZN(n682) );
NOR2_X1 U18272 ( .A1(n696), .A2(n697), .ZN(n690) );
NOR2_X1 U18273 ( .A1(n367), .A2(n692), .ZN(n691) );
NOR2_X1 U18274 ( .A1(n20005), .A2(n378), .ZN(n697) );
NAND2_X1 U18275 ( .A1(n652), .A2(n653), .ZN(n644) );
NOR2_X1 U18276 ( .A1(n658), .A2(n659), .ZN(n652) );
NOR2_X1 U18277 ( .A1(n367), .A2(n654), .ZN(n653) );
NOR2_X1 U18278 ( .A1(n20004), .A2(n378), .ZN(n659) );
NAND2_X1 U18279 ( .A1(n612), .A2(n613), .ZN(n604) );
NOR2_X1 U18280 ( .A1(n618), .A2(n619), .ZN(n612) );
NOR2_X1 U18281 ( .A1(n367), .A2(n614), .ZN(n613) );
NOR2_X1 U18282 ( .A1(n378), .A2(n20003), .ZN(n619) );
NAND2_X1 U18283 ( .A1(n572), .A2(n573), .ZN(n564) );
NOR2_X1 U18284 ( .A1(n578), .A2(n579), .ZN(n572) );
NOR2_X1 U18285 ( .A1(n367), .A2(n574), .ZN(n573) );
NOR2_X1 U18286 ( .A1(n20002), .A2(n378), .ZN(n579) );
NAND2_X1 U18287 ( .A1(n532), .A2(n533), .ZN(n524) );
NOR2_X1 U18288 ( .A1(n538), .A2(n539), .ZN(n532) );
NOR2_X1 U18289 ( .A1(n367), .A2(n534), .ZN(n533) );
NOR2_X1 U18290 ( .A1(n20001), .A2(n378), .ZN(n539) );
NOR2_X1 U18291 ( .A1(alu_operand_b_ex_4), .A2(n10005), .ZN(n10004) );
NOR2_X1 U18292 ( .A1(n10006), .A2(n10007), .ZN(n10005) );
NOR2_X1 U18293 ( .A1(n20864), .A2(n8115), .ZN(n10007) );
NOR2_X1 U18294 ( .A1(n9918), .A2(n10008), .ZN(n10006) );
NAND2_X1 U18295 ( .A1(n1426), .A2(n1427), .ZN(n32) );
NOR2_X1 U18296 ( .A1(n1430), .A2(n1431), .ZN(n1426) );
NOR2_X1 U18297 ( .A1(n20822), .A2(n20920), .ZN(n1427) );
NOR2_X1 U18298 ( .A1(n1432), .A2(n1433), .ZN(n1430) );
NOR2_X1 U18299 ( .A1(n883), .A2(n899), .ZN(n888) );
NAND2_X1 U18300 ( .A1(n16475), .A2(alu_operand_b_ex_1), .ZN(n899) );
NOR2_X1 U18301 ( .A1(n323), .A2(n337), .ZN(n328) );
NAND2_X1 U18302 ( .A1(n16474), .A2(alu_operand_b_ex_3), .ZN(n337) );
NOR2_X1 U18303 ( .A1(n282), .A2(n296), .ZN(n287) );
NAND2_X1 U18304 ( .A1(n16475), .A2(alu_operand_b_ex_4), .ZN(n296) );
NOR2_X1 U18305 ( .A1(n240), .A2(n254), .ZN(n245) );
NAND2_X1 U18306 ( .A1(n16474), .A2(n255), .ZN(n254) );
NOR2_X1 U18307 ( .A1(n16364), .A2(n20291), .ZN(n9091) );
NOR2_X1 U18308 ( .A1(n16364), .A2(n20330), .ZN(n9132) );
NOR2_X1 U18309 ( .A1(n16364), .A2(n20369), .ZN(n9173) );
NOR2_X1 U18310 ( .A1(n8601), .A2(n20408), .ZN(n9214) );
NOR2_X1 U18311 ( .A1(n8601), .A2(n20448), .ZN(n9255) );
NOR2_X1 U18312 ( .A1(n16364), .A2(n20252), .ZN(n9050) );
NAND2_X1 U18313 ( .A1(n1432), .A2(n9974), .ZN(n8430) );
NAND2_X1 U18314 ( .A1(n9975), .A2(n9976), .ZN(n9974) );
NOR2_X1 U18315 ( .A1(n10017), .A2(n10018), .ZN(n9975) );
NOR2_X1 U18316 ( .A1(n9977), .A2(n9978), .ZN(n9976) );
NOR2_X1 U18317 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
NAND2_X1 U18318 ( .A1(n16475), .A2(n1297), .ZN(n1296) );
NOR2_X1 U18319 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
NAND2_X1 U18320 ( .A1(n16474), .A2(n1219), .ZN(n1218) );
NOR2_X1 U18321 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND2_X1 U18322 ( .A1(n16474), .A2(n1180), .ZN(n1179) );
NOR2_X1 U18323 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NAND2_X1 U18324 ( .A1(n16474), .A2(n1141), .ZN(n1140) );
NOR2_X1 U18325 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND2_X1 U18326 ( .A1(n16474), .A2(n1005), .ZN(n1004) );
NOR2_X1 U18327 ( .A1(n965), .A2(n966), .ZN(n964) );
NAND2_X1 U18328 ( .A1(n16474), .A2(n967), .ZN(n966) );
NOR2_X1 U18329 ( .A1(n926), .A2(n927), .ZN(n925) );
NAND2_X1 U18330 ( .A1(n16475), .A2(n928), .ZN(n927) );
NOR2_X1 U18331 ( .A1(n845), .A2(n846), .ZN(n844) );
NAND2_X1 U18332 ( .A1(n16475), .A2(n847), .ZN(n846) );
NOR2_X1 U18333 ( .A1(n806), .A2(n807), .ZN(n805) );
NAND2_X1 U18334 ( .A1(n16475), .A2(n808), .ZN(n807) );
NOR2_X1 U18335 ( .A1(n768), .A2(n769), .ZN(n767) );
NAND2_X1 U18336 ( .A1(n16475), .A2(n770), .ZN(n769) );
NOR2_X1 U18337 ( .A1(n730), .A2(n731), .ZN(n729) );
NAND2_X1 U18338 ( .A1(n16475), .A2(n732), .ZN(n731) );
NOR2_X1 U18339 ( .A1(n693), .A2(n694), .ZN(n692) );
NAND2_X1 U18340 ( .A1(n16475), .A2(n695), .ZN(n694) );
NOR2_X1 U18341 ( .A1(n655), .A2(n656), .ZN(n654) );
NAND2_X1 U18342 ( .A1(n16475), .A2(n657), .ZN(n656) );
NOR2_X1 U18343 ( .A1(n615), .A2(n616), .ZN(n614) );
NAND2_X1 U18344 ( .A1(n16475), .A2(n617), .ZN(n616) );
NOR2_X1 U18345 ( .A1(n575), .A2(n576), .ZN(n574) );
NAND2_X1 U18346 ( .A1(n16475), .A2(n577), .ZN(n576) );
NOR2_X1 U18347 ( .A1(n535), .A2(n536), .ZN(n534) );
NAND2_X1 U18348 ( .A1(n16475), .A2(n537), .ZN(n536) );
NAND2_X1 U18349 ( .A1(n10315), .A2(n10316), .ZN(n3018) );
NOR2_X1 U18350 ( .A1(n10317), .A2(n10318), .ZN(n10316) );
NOR2_X1 U18351 ( .A1(n10321), .A2(n10322), .ZN(n10315) );
NAND2_X1 U18352 ( .A1(n5168), .A2(n5142), .ZN(n10318) );
NOR2_X1 U18353 ( .A1(n149), .A2(n169), .ZN(n156) );
NAND2_X1 U18354 ( .A1(n16475), .A2(n170), .ZN(n169) );
NOR2_X1 U18355 ( .A1(n20645), .A2(n971), .ZN(n968) );
NOR2_X1 U18356 ( .A1(n972), .A2(n973), .ZN(n971) );
NOR2_X1 U18357 ( .A1(n16476), .A2(n967), .ZN(n972) );
NAND2_X1 U18358 ( .A1(n974), .A2(n16473), .ZN(n973) );
NOR2_X1 U18359 ( .A1(n20329), .A2(n622), .ZN(n618) );
NOR2_X1 U18360 ( .A1(n623), .A2(n624), .ZN(n622) );
NOR2_X1 U18361 ( .A1(n15801), .A2(n617), .ZN(n623) );
NAND2_X1 U18362 ( .A1(n625), .A2(n16473), .ZN(n624) );
NOR2_X1 U18363 ( .A1(n16476), .A2(n465), .ZN(n456) );
NAND2_X1 U18364 ( .A1(n466), .A2(n20864), .ZN(n465) );
NOR2_X1 U18365 ( .A1(n15801), .A2(n211), .ZN(n202) );
NAND2_X1 U18366 ( .A1(n20841), .A2(n213), .ZN(n211) );
NOR2_X1 U18367 ( .A1(n20808), .A2(n1067), .ZN(n1063) );
NOR2_X1 U18368 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U18369 ( .A1(n16476), .A2(n1046), .ZN(n1068) );
NAND2_X1 U18370 ( .A1(n1070), .A2(n16473), .ZN(n1069) );
NOR2_X1 U18371 ( .A1(n20766), .A2(n419), .ZN(n415) );
NOR2_X1 U18372 ( .A1(n420), .A2(n421), .ZN(n419) );
NOR2_X1 U18373 ( .A1(n15801), .A2(n414), .ZN(n420) );
NAND2_X1 U18374 ( .A1(n422), .A2(n16473), .ZN(n421) );
NOR2_X1 U18375 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U18376 ( .A1(n16474), .A2(n1102), .ZN(n1101) );
NOR2_X1 U18377 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U18378 ( .A1(n16474), .A2(n1046), .ZN(n1045) );
NOR2_X1 U18379 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND2_X1 U18380 ( .A1(n16474), .A2(n1258), .ZN(n1257) );
NOR2_X1 U18381 ( .A1(n20845), .A2(n10009), .ZN(n10003) );
NOR2_X1 U18382 ( .A1(n10010), .A2(n10011), .ZN(n10009) );
NOR2_X1 U18383 ( .A1(n197), .A2(n8115), .ZN(n10011) );
NOR2_X1 U18384 ( .A1(n20827), .A2(n10012), .ZN(n10010) );
NOR2_X1 U18385 ( .A1(n20710), .A2(n1311), .ZN(n1309) );
NOR2_X1 U18386 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NOR2_X1 U18387 ( .A1(n1297), .A2(n15801), .ZN(n1312) );
NAND2_X1 U18388 ( .A1(n1314), .A2(n16473), .ZN(n1313) );
NOR2_X1 U18389 ( .A1(n20828), .A2(n1262), .ZN(n1260) );
NOR2_X1 U18390 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
NOR2_X1 U18391 ( .A1(n15801), .A2(n1258), .ZN(n1263) );
NAND2_X1 U18392 ( .A1(n1265), .A2(n16473), .ZN(n1264) );
NOR2_X1 U18393 ( .A1(n20702), .A2(n1223), .ZN(n1221) );
NOR2_X1 U18394 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NOR2_X1 U18395 ( .A1(n15801), .A2(n1219), .ZN(n1224) );
NAND2_X1 U18396 ( .A1(n1226), .A2(n16473), .ZN(n1225) );
NOR2_X1 U18397 ( .A1(n20698), .A2(n1184), .ZN(n1182) );
NOR2_X1 U18398 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NOR2_X1 U18399 ( .A1(n15801), .A2(n1180), .ZN(n1185) );
NAND2_X1 U18400 ( .A1(n1187), .A2(n16473), .ZN(n1186) );
NOR2_X1 U18401 ( .A1(n20694), .A2(n1145), .ZN(n1143) );
NOR2_X1 U18402 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NOR2_X1 U18403 ( .A1(n15801), .A2(n1141), .ZN(n1146) );
NAND2_X1 U18404 ( .A1(n1148), .A2(n16473), .ZN(n1147) );
NOR2_X1 U18405 ( .A1(n20679), .A2(n1009), .ZN(n1006) );
NOR2_X1 U18406 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NOR2_X1 U18407 ( .A1(n16476), .A2(n1005), .ZN(n1010) );
NAND2_X1 U18408 ( .A1(n1012), .A2(n16473), .ZN(n1011) );
NOR2_X1 U18409 ( .A1(n20607), .A2(n932), .ZN(n929) );
NOR2_X1 U18410 ( .A1(n933), .A2(n934), .ZN(n932) );
NOR2_X1 U18411 ( .A1(n16476), .A2(n928), .ZN(n933) );
NAND2_X1 U18412 ( .A1(n935), .A2(n16473), .ZN(n934) );
NOR2_X1 U18413 ( .A1(n20567), .A2(n851), .ZN(n848) );
NOR2_X1 U18414 ( .A1(n852), .A2(n853), .ZN(n851) );
NOR2_X1 U18415 ( .A1(n16476), .A2(n847), .ZN(n852) );
NAND2_X1 U18416 ( .A1(n854), .A2(n16473), .ZN(n853) );
NOR2_X1 U18417 ( .A1(n20527), .A2(n812), .ZN(n809) );
NOR2_X1 U18418 ( .A1(n813), .A2(n814), .ZN(n812) );
NOR2_X1 U18419 ( .A1(n15801), .A2(n808), .ZN(n813) );
NAND2_X1 U18420 ( .A1(n815), .A2(n16473), .ZN(n814) );
NOR2_X1 U18421 ( .A1(n20487), .A2(n774), .ZN(n771) );
NOR2_X1 U18422 ( .A1(n775), .A2(n776), .ZN(n774) );
NOR2_X1 U18423 ( .A1(n15801), .A2(n770), .ZN(n775) );
NAND2_X1 U18424 ( .A1(n777), .A2(n16473), .ZN(n776) );
NOR2_X1 U18425 ( .A1(n20447), .A2(n736), .ZN(n733) );
NOR2_X1 U18426 ( .A1(n737), .A2(n738), .ZN(n736) );
NOR2_X1 U18427 ( .A1(n16476), .A2(n732), .ZN(n737) );
NAND2_X1 U18428 ( .A1(n739), .A2(n16473), .ZN(n738) );
NOR2_X1 U18429 ( .A1(n20407), .A2(n699), .ZN(n696) );
NOR2_X1 U18430 ( .A1(n700), .A2(n701), .ZN(n699) );
NOR2_X1 U18431 ( .A1(n16476), .A2(n695), .ZN(n700) );
NAND2_X1 U18432 ( .A1(n702), .A2(n16473), .ZN(n701) );
NOR2_X1 U18433 ( .A1(n20368), .A2(n661), .ZN(n658) );
NOR2_X1 U18434 ( .A1(n662), .A2(n663), .ZN(n661) );
NOR2_X1 U18435 ( .A1(n15801), .A2(n657), .ZN(n662) );
NAND2_X1 U18436 ( .A1(n664), .A2(n16473), .ZN(n663) );
NOR2_X1 U18437 ( .A1(n20290), .A2(n582), .ZN(n578) );
NOR2_X1 U18438 ( .A1(n583), .A2(n584), .ZN(n582) );
NOR2_X1 U18439 ( .A1(n15801), .A2(n577), .ZN(n583) );
NAND2_X1 U18440 ( .A1(n585), .A2(n16473), .ZN(n584) );
NOR2_X1 U18441 ( .A1(n20251), .A2(n542), .ZN(n538) );
NOR2_X1 U18442 ( .A1(n543), .A2(n544), .ZN(n542) );
NOR2_X1 U18443 ( .A1(n16476), .A2(n537), .ZN(n543) );
NAND2_X1 U18444 ( .A1(n545), .A2(n16473), .ZN(n544) );
NOR2_X1 U18445 ( .A1(n20213), .A2(n502), .ZN(n498) );
NOR2_X1 U18446 ( .A1(n503), .A2(n504), .ZN(n502) );
NOR2_X1 U18447 ( .A1(n16476), .A2(n497), .ZN(n503) );
NAND2_X1 U18448 ( .A1(n505), .A2(n16473), .ZN(n504) );
NOR2_X1 U18449 ( .A1(n10013), .A2(n10014), .ZN(n10012) );
NAND2_X1 U18450 ( .A1(n20861), .A2(n20853), .ZN(n10014) );
NOR2_X1 U18451 ( .A1(n197), .A2(n10015), .ZN(n10013) );
NAND2_X1 U18452 ( .A1(n10016), .A2(alu_operand_b_ex_1), .ZN(n10015) );
NOR2_X1 U18453 ( .A1(n20718), .A2(n113), .ZN(n111) );
NOR2_X1 U18454 ( .A1(n114), .A2(n115), .ZN(n113) );
NOR2_X1 U18455 ( .A1(n16476), .A2(n109), .ZN(n114) );
NAND2_X1 U18456 ( .A1(n116), .A2(n16473), .ZN(n115) );
NOR2_X1 U18457 ( .A1(n20714), .A2(n58), .ZN(n56) );
NOR2_X1 U18458 ( .A1(n59), .A2(n60), .ZN(n58) );
NOR2_X1 U18459 ( .A1(n16476), .A2(n54), .ZN(n59) );
NAND2_X1 U18460 ( .A1(n61), .A2(n16473), .ZN(n60) );
NOR2_X1 U18461 ( .A1(n20810), .A2(n1106), .ZN(n1104) );
NOR2_X1 U18462 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR2_X1 U18463 ( .A1(n16476), .A2(n1102), .ZN(n1107) );
NAND2_X1 U18464 ( .A1(n1109), .A2(n16473), .ZN(n1108) );
NAND2_X1 U18465 ( .A1(n6265), .A2(n6266), .ZN(ex_block_i_alu_i_adder_in_a_26) );
NAND2_X1 U18466 ( .A1(n6238), .A2(n15870), .ZN(n6265) );
NAND2_X1 U18467 ( .A1(n16357), .A2(n655), .ZN(n6266) );
NAND2_X1 U18468 ( .A1(n6269), .A2(n6270), .ZN(ex_block_i_alu_i_adder_in_a_24) );
NAND2_X1 U18469 ( .A1(n6238), .A2(n15868), .ZN(n6269) );
NAND2_X1 U18470 ( .A1(n16357), .A2(n730), .ZN(n6270) );
NAND2_X1 U18471 ( .A1(n6267), .A2(n6268), .ZN(ex_block_i_alu_i_adder_in_a_25) );
NAND2_X1 U18472 ( .A1(n6238), .A2(n15869), .ZN(n6267) );
NAND2_X1 U18473 ( .A1(n16357), .A2(n693), .ZN(n6268) );
NAND2_X1 U18474 ( .A1(n6263), .A2(n6264), .ZN(ex_block_i_alu_i_adder_in_a_27) );
NAND2_X1 U18475 ( .A1(n16408), .A2(n15871), .ZN(n6263) );
NAND2_X1 U18476 ( .A1(n16357), .A2(n615), .ZN(n6264) );
NAND2_X1 U18477 ( .A1(n6261), .A2(n6262), .ZN(ex_block_i_alu_i_adder_in_a_28) );
NAND2_X1 U18478 ( .A1(n6238), .A2(n15872), .ZN(n6261) );
NAND2_X1 U18479 ( .A1(n16357), .A2(n575), .ZN(n6262) );
NAND2_X1 U18480 ( .A1(n6259), .A2(n6260), .ZN(ex_block_i_alu_i_adder_in_a_29) );
NAND2_X1 U18481 ( .A1(n16408), .A2(n15873), .ZN(n6259) );
NAND2_X1 U18482 ( .A1(n16357), .A2(n535), .ZN(n6260) );
NOR2_X1 U18483 ( .A1(n909), .A2(n910), .ZN(n907) );
NOR2_X1 U18484 ( .A1(n92), .A2(n20672), .ZN(n909) );
NOR2_X1 U18485 ( .A1(n90), .A2(n20753), .ZN(n910) );
NOR2_X1 U18486 ( .A1(n478), .A2(n479), .ZN(n476) );
NOR2_X1 U18487 ( .A1(n92), .A2(n20638), .ZN(n478) );
NOR2_X1 U18488 ( .A1(n16469), .A2(n20749), .ZN(n479) );
NOR2_X1 U18489 ( .A1(n348), .A2(n349), .ZN(n346) );
NOR2_X1 U18490 ( .A1(n92), .A2(n20584), .ZN(n348) );
NOR2_X1 U18491 ( .A1(n16469), .A2(n20743), .ZN(n349) );
NOR2_X1 U18492 ( .A1(n307), .A2(n308), .ZN(n305) );
NOR2_X1 U18493 ( .A1(n92), .A2(n20545), .ZN(n307) );
NOR2_X1 U18494 ( .A1(n16469), .A2(n20738), .ZN(n308) );
INV_X1 U18495 ( .A(n3412), .ZN(n20726) );
INV_X1 U18496 ( .A(n3407), .ZN(n20720) );
INV_X1 U18497 ( .A(n3402), .ZN(n19871) );
INV_X1 U18498 ( .A(n3397), .ZN(n19868) );
INV_X1 U18499 ( .A(n3553), .ZN(n19866) );
NAND2_X1 U18500 ( .A1(n16474), .A2(n54), .ZN(n52) );
NOR2_X1 U18501 ( .A1(n9990), .A2(n9991), .ZN(n9988) );
NOR2_X1 U18502 ( .A1(n9970), .A2(n1297), .ZN(n9991) );
NOR2_X1 U18503 ( .A1(n20864), .A2(n9992), .ZN(n9990) );
NOR2_X1 U18504 ( .A1(alu_operand_b_ex_1), .A2(n7571), .ZN(n9992) );
NAND2_X1 U18505 ( .A1(n492), .A2(n493), .ZN(n484) );
NOR2_X1 U18506 ( .A1(n367), .A2(n494), .ZN(n493) );
NOR2_X1 U18507 ( .A1(n498), .A2(n499), .ZN(n492) );
NOR2_X1 U18508 ( .A1(n495), .A2(n496), .ZN(n494) );
NAND2_X1 U18509 ( .A1(n6012), .A2(n6013), .ZN(ex_block_i_alu_i_adder_in_b_24) );
NOR2_X1 U18510 ( .A1(n6022), .A2(n6023), .ZN(n6012) );
NOR2_X1 U18511 ( .A1(n6014), .A2(n6015), .ZN(n6013) );
NOR2_X1 U18512 ( .A1(n5917), .A2(n16102), .ZN(n6022) );
NAND2_X1 U18513 ( .A1(n5970), .A2(n5971), .ZN(ex_block_i_alu_i_adder_in_b_27) );
NOR2_X1 U18514 ( .A1(n5980), .A2(n5981), .ZN(n5970) );
NOR2_X1 U18515 ( .A1(n5972), .A2(n5973), .ZN(n5971) );
NOR2_X1 U18516 ( .A1(n5917), .A2(n16099), .ZN(n5980) );
NAND2_X1 U18517 ( .A1(n5956), .A2(n5957), .ZN(ex_block_i_alu_i_adder_in_b_28) );
NOR2_X1 U18518 ( .A1(n5966), .A2(n5967), .ZN(n5956) );
NOR2_X1 U18519 ( .A1(n5958), .A2(n5959), .ZN(n5957) );
NOR2_X1 U18520 ( .A1(n5917), .A2(n16098), .ZN(n5966) );
NAND2_X1 U18521 ( .A1(n16472), .A2(n1297), .ZN(n1314) );
NAND2_X1 U18522 ( .A1(n16472), .A2(n109), .ZN(n116) );
NAND2_X1 U18523 ( .A1(n16472), .A2(n54), .ZN(n61) );
NAND2_X1 U18524 ( .A1(n16472), .A2(n808), .ZN(n815) );
NAND2_X1 U18525 ( .A1(n16472), .A2(n770), .ZN(n777) );
NAND2_X1 U18526 ( .A1(n16472), .A2(n732), .ZN(n739) );
NAND2_X1 U18527 ( .A1(n16472), .A2(n695), .ZN(n702) );
NAND2_X1 U18528 ( .A1(n16472), .A2(n657), .ZN(n664) );
NAND2_X1 U18529 ( .A1(n16472), .A2(n617), .ZN(n625) );
NAND2_X1 U18530 ( .A1(n16472), .A2(n577), .ZN(n585) );
NAND2_X1 U18531 ( .A1(n16472), .A2(n537), .ZN(n545) );
NAND2_X1 U18532 ( .A1(n16472), .A2(n497), .ZN(n505) );
NAND2_X1 U18533 ( .A1(n16472), .A2(n414), .ZN(n422) );
NAND2_X1 U18534 ( .A1(n16472), .A2(n1258), .ZN(n1265) );
NAND2_X1 U18535 ( .A1(n16472), .A2(n1219), .ZN(n1226) );
NAND2_X1 U18536 ( .A1(n16472), .A2(n1180), .ZN(n1187) );
NAND2_X1 U18537 ( .A1(n16472), .A2(n1141), .ZN(n1148) );
NAND2_X1 U18538 ( .A1(n16472), .A2(n1102), .ZN(n1109) );
NAND2_X1 U18539 ( .A1(n16472), .A2(n1046), .ZN(n1070) );
NAND2_X1 U18540 ( .A1(n16472), .A2(n1005), .ZN(n1012) );
NAND2_X1 U18541 ( .A1(n16472), .A2(n967), .ZN(n974) );
NAND2_X1 U18542 ( .A1(n16472), .A2(n928), .ZN(n935) );
NAND2_X1 U18543 ( .A1(n16472), .A2(n847), .ZN(n854) );
NAND2_X1 U18544 ( .A1(n3963), .A2(n3964), .ZN(n3548) );
NOR2_X1 U18545 ( .A1(n3777), .A2(n3970), .ZN(n3963) );
NOR2_X1 U18546 ( .A1(n3965), .A2(n3966), .ZN(n3964) );
NAND2_X1 U18547 ( .A1(n3971), .A2(n3972), .ZN(n3970) );
NAND2_X1 U18548 ( .A1(n5998), .A2(n5999), .ZN(ex_block_i_alu_i_adder_in_b_25) );
NOR2_X1 U18549 ( .A1(n6008), .A2(n6009), .ZN(n5998) );
NOR2_X1 U18550 ( .A1(n6000), .A2(n6001), .ZN(n5999) );
NOR2_X1 U18551 ( .A1(n5917), .A2(n16101), .ZN(n6008) );
NAND2_X1 U18552 ( .A1(n5984), .A2(n5985), .ZN(ex_block_i_alu_i_adder_in_b_26) );
NOR2_X1 U18553 ( .A1(n5994), .A2(n5995), .ZN(n5984) );
NOR2_X1 U18554 ( .A1(n5986), .A2(n5987), .ZN(n5985) );
NOR2_X1 U18555 ( .A1(n5917), .A2(n16100), .ZN(n5994) );
NAND2_X1 U18556 ( .A1(n5942), .A2(n5943), .ZN(ex_block_i_alu_i_adder_in_b_29) );
NOR2_X1 U18557 ( .A1(n5952), .A2(n5953), .ZN(n5942) );
NOR2_X1 U18558 ( .A1(n5944), .A2(n5945), .ZN(n5943) );
NOR2_X1 U18559 ( .A1(n5917), .A2(n16097), .ZN(n5952) );
NAND2_X1 U18560 ( .A1(n16474), .A2(n414), .ZN(n413) );
NAND2_X1 U18561 ( .A1(n16475), .A2(n109), .ZN(n108) );
NAND2_X1 U18562 ( .A1(n16475), .A2(n497), .ZN(n496) );
NAND2_X1 U18563 ( .A1(alu_operand_b_ex_2), .A2(n20871), .ZN(n10016) );
INV_X1 U18564 ( .A(n7693), .ZN(n20888) );
INV_X1 U18565 ( .A(n7654), .ZN(n20889) );
INV_X1 U18566 ( .A(instr_req_o), .ZN(n20879) );
NAND2_X1 U18567 ( .A1(n104), .A2(n105), .ZN(n96) );
NOR2_X1 U18568 ( .A1(n49), .A2(n106), .ZN(n105) );
NOR2_X1 U18569 ( .A1(n110), .A2(n111), .ZN(n104) );
NOR2_X1 U18570 ( .A1(n107), .A2(n108), .ZN(n106) );
NAND2_X1 U18571 ( .A1(n47), .A2(n48), .ZN(n36) );
NOR2_X1 U18572 ( .A1(n49), .A2(n50), .ZN(n48) );
NOR2_X1 U18573 ( .A1(n55), .A2(n56), .ZN(n47) );
NOR2_X1 U18574 ( .A1(n51), .A2(n52), .ZN(n50) );
NAND2_X1 U18575 ( .A1(n1292), .A2(n1293), .ZN(n1285) );
NOR2_X1 U18576 ( .A1(n1308), .A2(n1309), .ZN(n1292) );
NOR2_X1 U18577 ( .A1(n49), .A2(n1294), .ZN(n1293) );
NOR2_X1 U18578 ( .A1(n1320), .A2(n16335), .ZN(n1308) );
NAND2_X1 U18579 ( .A1(n1253), .A2(n1254), .ZN(n1246) );
NOR2_X1 U18580 ( .A1(n1259), .A2(n1260), .ZN(n1253) );
NOR2_X1 U18581 ( .A1(n49), .A2(n1255), .ZN(n1254) );
NOR2_X1 U18582 ( .A1(n1266), .A2(n16335), .ZN(n1259) );
NAND2_X1 U18583 ( .A1(n1214), .A2(n1215), .ZN(n1207) );
NOR2_X1 U18584 ( .A1(n1220), .A2(n1221), .ZN(n1214) );
NOR2_X1 U18585 ( .A1(n49), .A2(n1216), .ZN(n1215) );
NOR2_X1 U18586 ( .A1(n1227), .A2(n16335), .ZN(n1220) );
NAND2_X1 U18587 ( .A1(n1175), .A2(n1176), .ZN(n1168) );
NOR2_X1 U18588 ( .A1(n1181), .A2(n1182), .ZN(n1175) );
NOR2_X1 U18589 ( .A1(n49), .A2(n1177), .ZN(n1176) );
NOR2_X1 U18590 ( .A1(n1188), .A2(n33), .ZN(n1181) );
NAND2_X1 U18591 ( .A1(n1136), .A2(n1137), .ZN(n1129) );
NOR2_X1 U18592 ( .A1(n1142), .A2(n1143), .ZN(n1136) );
NOR2_X1 U18593 ( .A1(n49), .A2(n1138), .ZN(n1137) );
NOR2_X1 U18594 ( .A1(n1149), .A2(n16335), .ZN(n1142) );
NAND2_X1 U18595 ( .A1(n1097), .A2(n1098), .ZN(n1090) );
NOR2_X1 U18596 ( .A1(n1103), .A2(n1104), .ZN(n1097) );
NOR2_X1 U18597 ( .A1(n49), .A2(n1099), .ZN(n1098) );
NOR2_X1 U18598 ( .A1(n1110), .A2(n33), .ZN(n1103) );
NAND2_X1 U18599 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
NAND2_X1 U18600 ( .A1(n16471), .A2(n1331), .ZN(n1330) );
NOR2_X1 U18601 ( .A1(n1332), .A2(n1333), .ZN(n1329) );
NOR2_X1 U18602 ( .A1(n16470), .A2(n16232), .ZN(n1332) );
NAND2_X1 U18603 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U18604 ( .A1(n16471), .A2(n1275), .ZN(n1274) );
NOR2_X1 U18605 ( .A1(n1276), .A2(n1277), .ZN(n1273) );
NOR2_X1 U18606 ( .A1(n16470), .A2(n16214), .ZN(n1276) );
NAND2_X1 U18607 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND2_X1 U18608 ( .A1(n16471), .A2(n1236), .ZN(n1235) );
NOR2_X1 U18609 ( .A1(n1237), .A2(n1238), .ZN(n1234) );
NOR2_X1 U18610 ( .A1(n16470), .A2(n16211), .ZN(n1237) );
NAND2_X1 U18611 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NAND2_X1 U18612 ( .A1(n16471), .A2(n1197), .ZN(n1196) );
NOR2_X1 U18613 ( .A1(n1198), .A2(n1199), .ZN(n1195) );
NOR2_X1 U18614 ( .A1(n16470), .A2(n16229), .ZN(n1198) );
NAND2_X1 U18615 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U18616 ( .A1(n16471), .A2(n1158), .ZN(n1157) );
NOR2_X1 U18617 ( .A1(n1159), .A2(n1160), .ZN(n1156) );
NOR2_X1 U18618 ( .A1(n16470), .A2(n16226), .ZN(n1159) );
NAND2_X1 U18619 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U18620 ( .A1(n16471), .A2(n1119), .ZN(n1118) );
NOR2_X1 U18621 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
NOR2_X1 U18622 ( .A1(n16470), .A2(n16223), .ZN(n1120) );
AND2_X1 U18623 ( .A1(n10348), .A2(n7653), .ZN(n7622) );
NOR2_X1 U18624 ( .A1(n20888), .A2(n20889), .ZN(n10348) );
NAND2_X1 U18625 ( .A1(n3967), .A2(n3968), .ZN(n3966) );
NAND2_X1 U18626 ( .A1(n3774), .A2(crash_dump_o_11_), .ZN(n3967) );
NAND2_X1 U18627 ( .A1(n3773), .A2(data_addr_o_11_), .ZN(n3968) );
NAND2_X1 U18628 ( .A1(n1041), .A2(n1042), .ZN(n1031) );
NOR2_X1 U18629 ( .A1(n1063), .A2(n1064), .ZN(n1041) );
NOR2_X1 U18630 ( .A1(n367), .A2(n1043), .ZN(n1042) );
NOR2_X1 U18631 ( .A1(n20013), .A2(n378), .ZN(n1064) );
NAND2_X1 U18632 ( .A1(n1000), .A2(n1001), .ZN(n993) );
NOR2_X1 U18633 ( .A1(n1006), .A2(n1007), .ZN(n1000) );
NOR2_X1 U18634 ( .A1(n367), .A2(n1002), .ZN(n1001) );
NOR2_X1 U18635 ( .A1(n20012), .A2(n378), .ZN(n1007) );
NAND2_X1 U18636 ( .A1(n962), .A2(n963), .ZN(n954) );
NOR2_X1 U18637 ( .A1(n968), .A2(n969), .ZN(n962) );
NOR2_X1 U18638 ( .A1(n367), .A2(n964), .ZN(n963) );
NOR2_X1 U18639 ( .A1(n378), .A2(n20011), .ZN(n969) );
NAND2_X1 U18640 ( .A1(n409), .A2(n410), .ZN(n401) );
NOR2_X1 U18641 ( .A1(n367), .A2(n411), .ZN(n410) );
NOR2_X1 U18642 ( .A1(n415), .A2(n416), .ZN(n409) );
NOR2_X1 U18643 ( .A1(n412), .A2(n413), .ZN(n411) );
NAND2_X1 U18644 ( .A1(n902), .A2(n903), .ZN(n901) );
NAND2_X1 U18645 ( .A1(n16471), .A2(n904), .ZN(n903) );
NOR2_X1 U18646 ( .A1(n905), .A2(n906), .ZN(n902) );
NOR2_X1 U18647 ( .A1(n83), .A2(n16208), .ZN(n905) );
NAND2_X1 U18648 ( .A1(n470), .A2(n471), .ZN(n469) );
NAND2_X1 U18649 ( .A1(n78), .A2(n472), .ZN(n471) );
NOR2_X1 U18650 ( .A1(n473), .A2(n474), .ZN(n470) );
NOR2_X1 U18651 ( .A1(n16470), .A2(n16205), .ZN(n473) );
NAND2_X1 U18652 ( .A1(n340), .A2(n341), .ZN(n339) );
NAND2_X1 U18653 ( .A1(n78), .A2(n342), .ZN(n341) );
NOR2_X1 U18654 ( .A1(n343), .A2(n344), .ZN(n340) );
NOR2_X1 U18655 ( .A1(n83), .A2(n16202), .ZN(n343) );
NAND2_X1 U18656 ( .A1(n299), .A2(n300), .ZN(n298) );
NAND2_X1 U18657 ( .A1(n78), .A2(n301), .ZN(n300) );
NOR2_X1 U18658 ( .A1(n302), .A2(n303), .ZN(n299) );
NOR2_X1 U18659 ( .A1(n83), .A2(n16244), .ZN(n302) );
NAND2_X1 U18660 ( .A1(n216), .A2(n217), .ZN(n215) );
NAND2_X1 U18661 ( .A1(n78), .A2(n218), .ZN(n217) );
NOR2_X1 U18662 ( .A1(n219), .A2(n220), .ZN(n216) );
NOR2_X1 U18663 ( .A1(n83), .A2(n16238), .ZN(n219) );
NAND2_X1 U18664 ( .A1(n173), .A2(n174), .ZN(n172) );
NAND2_X1 U18665 ( .A1(n78), .A2(n175), .ZN(n174) );
NOR2_X1 U18666 ( .A1(n176), .A2(n177), .ZN(n173) );
NOR2_X1 U18667 ( .A1(n83), .A2(n16220), .ZN(n176) );
NAND2_X1 U18668 ( .A1(n125), .A2(n126), .ZN(n124) );
NAND2_X1 U18669 ( .A1(n78), .A2(n127), .ZN(n126) );
NOR2_X1 U18670 ( .A1(n128), .A2(n129), .ZN(n125) );
NOR2_X1 U18671 ( .A1(n83), .A2(n16217), .ZN(n128) );
NAND2_X1 U18672 ( .A1(n76), .A2(n77), .ZN(n75) );
NAND2_X1 U18673 ( .A1(n78), .A2(n79), .ZN(n77) );
NOR2_X1 U18674 ( .A1(n80), .A2(n81), .ZN(n76) );
NOR2_X1 U18675 ( .A1(n83), .A2(n16235), .ZN(n80) );
NAND2_X1 U18676 ( .A1(n6002), .A2(n6003), .ZN(n6001) );
NAND2_X1 U18677 ( .A1(n695), .A2(n16334), .ZN(n6002) );
NAND2_X1 U18678 ( .A1(n20784), .A2(n5826), .ZN(n6003) );
INV_X1 U18679 ( .A(n695), .ZN(n20784) );
NAND2_X1 U18680 ( .A1(n5988), .A2(n5989), .ZN(n5987) );
NAND2_X1 U18681 ( .A1(n657), .A2(n16334), .ZN(n5988) );
NAND2_X1 U18682 ( .A1(n20781), .A2(n16409), .ZN(n5989) );
INV_X1 U18683 ( .A(n657), .ZN(n20781) );
NAND2_X1 U18684 ( .A1(n5974), .A2(n5975), .ZN(n5973) );
NAND2_X1 U18685 ( .A1(n617), .A2(n5904), .ZN(n5974) );
NAND2_X1 U18686 ( .A1(n20778), .A2(n5826), .ZN(n5975) );
INV_X1 U18687 ( .A(n617), .ZN(n20778) );
NAND2_X1 U18688 ( .A1(n5960), .A2(n5961), .ZN(n5959) );
NAND2_X1 U18689 ( .A1(n577), .A2(n16334), .ZN(n5960) );
NAND2_X1 U18690 ( .A1(n20775), .A2(n16409), .ZN(n5961) );
INV_X1 U18691 ( .A(n577), .ZN(n20775) );
NAND2_X1 U18692 ( .A1(n5946), .A2(n5947), .ZN(n5945) );
NAND2_X1 U18693 ( .A1(n537), .A2(n5904), .ZN(n5946) );
NAND2_X1 U18694 ( .A1(n20772), .A2(n5826), .ZN(n5947) );
INV_X1 U18695 ( .A(n537), .ZN(n20772) );
NAND2_X1 U18696 ( .A1(n6016), .A2(n6017), .ZN(n6015) );
NAND2_X1 U18697 ( .A1(n732), .A2(n16334), .ZN(n6016) );
NAND2_X1 U18698 ( .A1(n20787), .A2(n16409), .ZN(n6017) );
INV_X1 U18699 ( .A(n732), .ZN(n20787) );
NAND2_X1 U18700 ( .A1(n449), .A2(n450), .ZN(n442) );
NOR2_X1 U18701 ( .A1(n456), .A2(n457), .ZN(n449) );
NAND2_X1 U18702 ( .A1(n451), .A2(alu_operand_b_ex_2), .ZN(n450) );
NOR2_X1 U18703 ( .A1(n458), .A2(n33), .ZN(n457) );
NAND2_X1 U18704 ( .A1(n237), .A2(n238), .ZN(n230) );
NOR2_X1 U18705 ( .A1(n245), .A2(n246), .ZN(n237) );
NAND2_X1 U18706 ( .A1(n239), .A2(n240), .ZN(n238) );
NOR2_X1 U18707 ( .A1(n247), .A2(n16335), .ZN(n246) );
NAND2_X1 U18708 ( .A1(n5142), .A2(n20879), .ZN(n10302) );
NAND2_X1 U18709 ( .A1(n194), .A2(n195), .ZN(n187) );
NOR2_X1 U18710 ( .A1(n202), .A2(n203), .ZN(n194) );
NAND2_X1 U18711 ( .A1(n196), .A2(n197), .ZN(n195) );
NOR2_X1 U18712 ( .A1(n204), .A2(n33), .ZN(n203) );
NAND2_X1 U18713 ( .A1(n146), .A2(n147), .ZN(n139) );
NOR2_X1 U18714 ( .A1(n156), .A2(n157), .ZN(n146) );
NAND2_X1 U18715 ( .A1(n148), .A2(n149), .ZN(n147) );
NOR2_X1 U18716 ( .A1(n158), .A2(n16335), .ZN(n157) );
NAND2_X1 U18717 ( .A1(n871), .A2(n872), .ZN(rf_wdata_wb_ecc_o_1_) );
NOR2_X1 U18718 ( .A1(n900), .A2(n901), .ZN(n871) );
NOR2_X1 U18719 ( .A1(n873), .A2(n874), .ZN(n872) );
NAND2_X1 U18720 ( .A1(n907), .A2(n908), .ZN(n900) );
NAND2_X1 U18721 ( .A1(n440), .A2(n441), .ZN(rf_wdata_wb_ecc_o_2_) );
NOR2_X1 U18722 ( .A1(n468), .A2(n469), .ZN(n440) );
NOR2_X1 U18723 ( .A1(n442), .A2(n443), .ZN(n441) );
NAND2_X1 U18724 ( .A1(n476), .A2(n477), .ZN(n468) );
NAND2_X1 U18725 ( .A1(n311), .A2(n312), .ZN(rf_wdata_wb_ecc_o_3_) );
NOR2_X1 U18726 ( .A1(n338), .A2(n339), .ZN(n311) );
NOR2_X1 U18727 ( .A1(n313), .A2(n314), .ZN(n312) );
NAND2_X1 U18728 ( .A1(n346), .A2(n347), .ZN(n338) );
NAND2_X1 U18729 ( .A1(n270), .A2(n271), .ZN(rf_wdata_wb_ecc_o_4_) );
NOR2_X1 U18730 ( .A1(n297), .A2(n298), .ZN(n270) );
NOR2_X1 U18731 ( .A1(n272), .A2(n273), .ZN(n271) );
NAND2_X1 U18732 ( .A1(n305), .A2(n306), .ZN(n297) );
NAND2_X1 U18733 ( .A1(n228), .A2(n229), .ZN(rf_wdata_wb_ecc_o_5_) );
NOR2_X1 U18734 ( .A1(n256), .A2(n257), .ZN(n228) );
NOR2_X1 U18735 ( .A1(n230), .A2(n231), .ZN(n229) );
NAND2_X1 U18736 ( .A1(n258), .A2(n259), .ZN(n257) );
NAND2_X1 U18737 ( .A1(n185), .A2(n186), .ZN(rf_wdata_wb_ecc_o_6_) );
NOR2_X1 U18738 ( .A1(n187), .A2(n188), .ZN(n186) );
NOR2_X1 U18739 ( .A1(n214), .A2(n215), .ZN(n185) );
NAND2_X1 U18740 ( .A1(n189), .A2(n190), .ZN(n188) );
NAND2_X1 U18741 ( .A1(n137), .A2(n138), .ZN(rf_wdata_wb_ecc_o_7_) );
NOR2_X1 U18742 ( .A1(n139), .A2(n140), .ZN(n138) );
NOR2_X1 U18743 ( .A1(n171), .A2(n172), .ZN(n137) );
NAND2_X1 U18744 ( .A1(n141), .A2(n142), .ZN(n140) );
NAND2_X1 U18745 ( .A1(n94), .A2(n95), .ZN(rf_wdata_wb_ecc_o_8_) );
NOR2_X1 U18746 ( .A1(n96), .A2(n97), .ZN(n95) );
NOR2_X1 U18747 ( .A1(n123), .A2(n124), .ZN(n94) );
NAND2_X1 U18748 ( .A1(n98), .A2(n99), .ZN(n97) );
NAND2_X1 U18749 ( .A1(n10300), .A2(n10301), .ZN(core_busy_o) );
NOR2_X1 U18750 ( .A1(n10462), .A2(n10463), .ZN(n10300) );
NOR2_X1 U18751 ( .A1(n10302), .A2(n10303), .ZN(n10301) );
OR2_X1 U18752 ( .A1(n3704), .A2(n15878), .ZN(n10463) );
NAND2_X1 U18753 ( .A1(n20990), .A2(alu_operand_b_ex_4), .ZN(n5801) );
NAND2_X1 U18754 ( .A1(ex_block_i_alu_i_shift_amt_compl_4), .A2(n1444), .ZN(n5800) );
NOR2_X1 U18755 ( .A1(n21661), .A2(n21660), .ZN(ex_block_i_alu_i_shift_amt_compl_4) );
BUF_X1 U18756 ( .A(n1706), .Z(n16459) );
NAND2_X1 U18757 ( .A1(n5954), .A2(n5955), .ZN(n5953) );
NAND2_X1 U18758 ( .A1(n16410), .A2(n20252), .ZN(n5955) );
NAND2_X1 U18759 ( .A1(n5916), .A2(n20773), .ZN(n5954) );
NAND2_X1 U18760 ( .A1(n5930), .A2(n5931), .ZN(n5929) );
NAND2_X1 U18761 ( .A1(n5818), .A2(n20214), .ZN(n5931) );
NAND2_X1 U18762 ( .A1(n5916), .A2(n20770), .ZN(n5930) );
NAND2_X1 U18763 ( .A1(n5914), .A2(n5915), .ZN(n5913) );
NAND2_X1 U18764 ( .A1(n16410), .A2(n20176), .ZN(n5915) );
NAND2_X1 U18765 ( .A1(n5916), .A2(n20767), .ZN(n5914) );
NOR2_X1 U18766 ( .A1(n10344), .A2(n7629), .ZN(n7684) );
NAND2_X1 U18767 ( .A1(n7620), .A2(n7700), .ZN(n10344) );
NAND2_X1 U18768 ( .A1(n5805), .A2(n5806), .ZN(ex_block_i_alu_i_shift_amt_2) );
NAND2_X1 U18769 ( .A1(n20990), .A2(alu_operand_b_ex_2), .ZN(n5806) );
NAND2_X1 U18770 ( .A1(ex_block_i_alu_i_shift_amt_compl_2), .A2(n1444), .ZN(n5805) );
NOR2_X1 U18771 ( .A1(n21652), .A2(n21651), .ZN(ex_block_i_alu_i_shift_amt_compl_2) );
NOR2_X1 U18772 ( .A1(alu_operand_b_ex_3), .A2(n20864), .ZN(n9944) );
NOR2_X1 U18773 ( .A1(n7646), .A2(n7643), .ZN(n7678) );
NOR2_X1 U18774 ( .A1(n359), .A2(n20681), .ZN(n1081) );
NOR2_X1 U18775 ( .A1(n359), .A2(n20672), .ZN(n1023) );
NOR2_X1 U18776 ( .A1(n359), .A2(n20638), .ZN(n985) );
NAND2_X1 U18777 ( .A1(n9917), .A2(n7719), .ZN(n8312) );
NOR2_X1 U18778 ( .A1(alu_operand_b_ex_4), .A2(n9918), .ZN(n9917) );
NAND2_X1 U18779 ( .A1(n5807), .A2(n5808), .ZN(ex_block_i_alu_i_shift_amt_1) );
NAND2_X1 U18780 ( .A1(n20990), .A2(alu_operand_b_ex_1), .ZN(n5808) );
NAND2_X1 U18781 ( .A1(ex_block_i_alu_i_shift_amt_compl_1), .A2(n1444), .ZN(n5807) );
NAND2_X1 U18782 ( .A1(n21650), .A2(n21649), .ZN(ex_block_i_alu_i_shift_amt_compl_1) );
NAND2_X1 U18783 ( .A1(n5803), .A2(n5804), .ZN(ex_block_i_alu_i_shift_amt_3) );
NAND2_X1 U18784 ( .A1(n20990), .A2(alu_operand_b_ex_3), .ZN(n5804) );
NAND2_X1 U18785 ( .A1(ex_block_i_alu_i_shift_amt_compl_3), .A2(n1444), .ZN(n5803) );
NOR2_X1 U18786 ( .A1(n21656), .A2(n21655), .ZN(ex_block_i_alu_i_shift_amt_compl_3) );
NOR2_X1 U18787 ( .A1(n7699), .A2(n7700), .ZN(n7619) );
NAND2_X1 U18788 ( .A1(n7658), .A2(n20885), .ZN(n7699) );
NOR2_X1 U18789 ( .A1(n20584), .A2(n359), .ZN(n946) );
NOR2_X1 U18790 ( .A1(n20545), .A2(n359), .ZN(n865) );
NAND2_X1 U18791 ( .A1(n10128), .A2(n10129), .ZN(n10115) );
NAND2_X1 U18792 ( .A1(n20761), .A2(n5799), .ZN(n10128) );
NAND2_X1 U18793 ( .A1(n20136), .A2(n10130), .ZN(n10129) );
NAND2_X1 U18794 ( .A1(n16467), .A2(n693), .ZN(n5741) );
NAND2_X1 U18795 ( .A1(n16466), .A2(n170), .ZN(n5742) );
NAND2_X1 U18796 ( .A1(n16467), .A2(n730), .ZN(n5739) );
NAND2_X1 U18797 ( .A1(n16466), .A2(n107), .ZN(n5740) );
NAND2_X1 U18798 ( .A1(n5809), .A2(n5810), .ZN(ex_block_i_alu_i_shift_amt_0) );
NAND2_X1 U18799 ( .A1(ex_block_i_alu_i_shift_amt_compl_0), .A2(n1444), .ZN(n5809) );
NAND2_X1 U18800 ( .A1(n20990), .A2(ex_block_i_alu_i_shift_amt_compl_0), .ZN(n5810) );
NAND2_X1 U18801 ( .A1(n16467), .A2(n1217), .ZN(n5777) );
NAND2_X1 U18802 ( .A1(n1338), .A2(n926), .ZN(n5778) );
NAND2_X1 U18803 ( .A1(n16468), .A2(n1102), .ZN(n5783) );
NAND2_X1 U18804 ( .A1(n1338), .A2(n1046), .ZN(n5784) );
NAND2_X1 U18805 ( .A1(n16468), .A2(n1295), .ZN(n5771) );
NAND2_X1 U18806 ( .A1(n1338), .A2(n806), .ZN(n5772) );
NAND2_X1 U18807 ( .A1(n1338), .A2(n1391), .ZN(n5798) );
INV_X1 U18808 ( .A(n10130), .ZN(n20761) );
NOR2_X1 U18809 ( .A1(n8601), .A2(n20137), .ZN(n10135) );
NOR2_X1 U18810 ( .A1(alu_operand_b_ex_2), .A2(n21653), .ZN(n21651) );
NOR2_X1 U18811 ( .A1(alu_operand_b_ex_3), .A2(n21654), .ZN(n21655) );
NOR2_X1 U18812 ( .A1(alu_operand_b_ex_4), .A2(n21659), .ZN(n21660) );
NOR2_X1 U18813 ( .A1(n16405), .A2(n6525), .ZN(n6524) );
NOR2_X1 U18814 ( .A1(n16364), .A2(n20176), .ZN(n8964) );
NOR2_X1 U18815 ( .A1(n16364), .A2(n20214), .ZN(n9009) );
NOR2_X1 U18816 ( .A1(n20872), .A2(n16462), .ZN(n6503) );
NOR2_X1 U18817 ( .A1(n20870), .A2(n1566), .ZN(n6437) );
NOR2_X1 U18818 ( .A1(n20831), .A2(n16462), .ZN(n6497) );
NOR2_X1 U18819 ( .A1(n20829), .A2(n16462), .ZN(n6491) );
NOR2_X1 U18820 ( .A1(n20817), .A2(n16462), .ZN(n6485) );
NOR2_X1 U18821 ( .A1(n20815), .A2(n16462), .ZN(n6479) );
NOR2_X1 U18822 ( .A1(n20813), .A2(n16462), .ZN(n6473) );
NOR2_X1 U18823 ( .A1(n20811), .A2(n16462), .ZN(n6467) );
NOR2_X1 U18824 ( .A1(n20809), .A2(n16462), .ZN(n6461) );
NOR2_X1 U18825 ( .A1(n20806), .A2(n16462), .ZN(n6455) );
NOR2_X1 U18826 ( .A1(n20803), .A2(n16462), .ZN(n6449) );
NOR2_X1 U18827 ( .A1(n20800), .A2(n16462), .ZN(n6443) );
NOR2_X1 U18828 ( .A1(n20797), .A2(n1566), .ZN(n6431) );
NOR2_X1 U18829 ( .A1(n20794), .A2(n1566), .ZN(n6425) );
NOR2_X1 U18830 ( .A1(n20791), .A2(n1566), .ZN(n6419) );
NOR2_X1 U18831 ( .A1(n20788), .A2(n1566), .ZN(n6413) );
NOR2_X1 U18832 ( .A1(n20785), .A2(n1566), .ZN(n6407) );
NOR2_X1 U18833 ( .A1(n20782), .A2(n1566), .ZN(n6401) );
NOR2_X1 U18834 ( .A1(n20779), .A2(n1566), .ZN(n6395) );
NOR2_X1 U18835 ( .A1(n20776), .A2(n1566), .ZN(n6389) );
NOR2_X1 U18836 ( .A1(n20773), .A2(n1566), .ZN(n6383) );
NOR2_X1 U18837 ( .A1(n20770), .A2(n1566), .ZN(n6377) );
NOR2_X1 U18838 ( .A1(n20806), .A2(n16407), .ZN(n6436) );
NOR2_X1 U18839 ( .A1(n20803), .A2(n16406), .ZN(n6370) );
NOR2_X1 U18840 ( .A1(n20800), .A2(n16406), .ZN(n6352) );
NOR2_X1 U18841 ( .A1(n20797), .A2(n16406), .ZN(n6346) );
NOR2_X1 U18842 ( .A1(n20794), .A2(n16406), .ZN(n6340) );
NOR2_X1 U18843 ( .A1(n20791), .A2(n16406), .ZN(n6334) );
NOR2_X1 U18844 ( .A1(n20788), .A2(n16406), .ZN(n6328) );
NOR2_X1 U18845 ( .A1(n20785), .A2(n16406), .ZN(n6322) );
NOR2_X1 U18846 ( .A1(n20782), .A2(n16406), .ZN(n6314) );
NOR2_X1 U18847 ( .A1(n20870), .A2(n16407), .ZN(n6454) );
NOR2_X1 U18848 ( .A1(n20865), .A2(n16407), .ZN(n6448) );
NOR2_X1 U18849 ( .A1(n20862), .A2(n16407), .ZN(n6442) );
NOR2_X1 U18850 ( .A1(n20854), .A2(n16407), .ZN(n6430) );
NOR2_X1 U18851 ( .A1(n20847), .A2(n16407), .ZN(n6424) );
NOR2_X1 U18852 ( .A1(n20842), .A2(n16407), .ZN(n6418) );
NOR2_X1 U18853 ( .A1(n20840), .A2(n16407), .ZN(n6412) );
NOR2_X1 U18854 ( .A1(n20836), .A2(n16407), .ZN(n6406) );
NOR2_X1 U18855 ( .A1(n20834), .A2(n16407), .ZN(n6400) );
NOR2_X1 U18856 ( .A1(n20831), .A2(n16407), .ZN(n6394) );
NOR2_X1 U18857 ( .A1(n20829), .A2(n16407), .ZN(n6388) );
NOR2_X1 U18858 ( .A1(n20817), .A2(n16406), .ZN(n6382) );
NOR2_X1 U18859 ( .A1(n20815), .A2(n16406), .ZN(n6376) );
NOR2_X1 U18860 ( .A1(n20813), .A2(n16406), .ZN(n6364) );
NOR2_X1 U18861 ( .A1(n20811), .A2(n16406), .ZN(n6358) );
NOR2_X1 U18862 ( .A1(n20782), .A2(n6318), .ZN(n6438) );
NOR2_X1 U18863 ( .A1(n20831), .A2(n6318), .ZN(n6450) );
NOR2_X1 U18864 ( .A1(n20829), .A2(n6318), .ZN(n6444) );
NOR2_X1 U18865 ( .A1(n20817), .A2(n6318), .ZN(n6432) );
NOR2_X1 U18866 ( .A1(n20815), .A2(n6318), .ZN(n6426) );
NOR2_X1 U18867 ( .A1(n20813), .A2(n6318), .ZN(n6420) );
NOR2_X1 U18868 ( .A1(n20811), .A2(n6318), .ZN(n6414) );
NOR2_X1 U18869 ( .A1(n20809), .A2(n6318), .ZN(n6408) );
NOR2_X1 U18870 ( .A1(n20806), .A2(n6318), .ZN(n6402) );
NOR2_X1 U18871 ( .A1(n20803), .A2(n6318), .ZN(n6396) );
NOR2_X1 U18872 ( .A1(n20800), .A2(n6318), .ZN(n6390) );
NOR2_X1 U18873 ( .A1(n20785), .A2(n16405), .ZN(n6504) );
NOR2_X1 U18874 ( .A1(n20870), .A2(n16405), .ZN(n6317) );
NOR2_X1 U18875 ( .A1(n20865), .A2(n16405), .ZN(n6498) );
NOR2_X1 U18876 ( .A1(n20862), .A2(n16405), .ZN(n6492) );
NOR2_X1 U18877 ( .A1(n20854), .A2(n16405), .ZN(n6486) );
NOR2_X1 U18878 ( .A1(n20847), .A2(n16405), .ZN(n6480) );
NOR2_X1 U18879 ( .A1(n20842), .A2(n16405), .ZN(n6474) );
NOR2_X1 U18880 ( .A1(n20840), .A2(n16405), .ZN(n6468) );
NOR2_X1 U18881 ( .A1(n20836), .A2(n16405), .ZN(n6462) );
NOR2_X1 U18882 ( .A1(n20834), .A2(n16405), .ZN(n6456) );
NOR2_X1 U18883 ( .A1(n20865), .A2(n1566), .ZN(n6371) );
NOR2_X1 U18884 ( .A1(n20862), .A2(n1566), .ZN(n6353) );
NOR2_X1 U18885 ( .A1(n20854), .A2(n1566), .ZN(n6347) );
NOR2_X1 U18886 ( .A1(n20847), .A2(n1566), .ZN(n6341) );
NOR2_X1 U18887 ( .A1(n20842), .A2(n1566), .ZN(n6335) );
NOR2_X1 U18888 ( .A1(n20840), .A2(n1566), .ZN(n6329) );
NOR2_X1 U18889 ( .A1(n20836), .A2(n1566), .ZN(n6323) );
NOR2_X1 U18890 ( .A1(n20834), .A2(n1566), .ZN(n6316) );
NOR2_X1 U18891 ( .A1(n20767), .A2(n1566), .ZN(n6365) );
NOR2_X1 U18892 ( .A1(n20764), .A2(n1566), .ZN(n6359) );
NOR2_X1 U18893 ( .A1(n20779), .A2(n16405), .ZN(n6372) );
NOR2_X1 U18894 ( .A1(n20776), .A2(n16405), .ZN(n6354) );
NOR2_X1 U18895 ( .A1(n20773), .A2(n16405), .ZN(n6348) );
NOR2_X1 U18896 ( .A1(n20770), .A2(n16405), .ZN(n6342) );
NOR2_X1 U18897 ( .A1(n20767), .A2(n16405), .ZN(n6336) );
NOR2_X1 U18898 ( .A1(n20764), .A2(n16405), .ZN(n6330) );
NOR2_X1 U18899 ( .A1(n20872), .A2(n16405), .ZN(n6324) );
NOR2_X1 U18900 ( .A1(n20797), .A2(n16405), .ZN(n6384) );
NOR2_X1 U18901 ( .A1(n20794), .A2(n6318), .ZN(n6378) );
NOR2_X1 U18902 ( .A1(n20791), .A2(n6318), .ZN(n6366) );
NOR2_X1 U18903 ( .A1(n20788), .A2(n6318), .ZN(n6360) );
INV_X1 U18904 ( .A(n5799), .ZN(n20136) );
NOR2_X1 U18905 ( .A1(n20809), .A2(n16407), .ZN(n6502) );
NOR2_X1 U18906 ( .A1(n20779), .A2(n16406), .ZN(n6496) );
NOR2_X1 U18907 ( .A1(n20776), .A2(n16407), .ZN(n6490) );
NOR2_X1 U18908 ( .A1(n20773), .A2(n16406), .ZN(n6484) );
NOR2_X1 U18909 ( .A1(n20770), .A2(n16407), .ZN(n6478) );
NOR2_X1 U18910 ( .A1(n20767), .A2(n16406), .ZN(n6472) );
NOR2_X1 U18911 ( .A1(n20764), .A2(n16407), .ZN(n6466) );
NOR2_X1 U18912 ( .A1(n20872), .A2(n16406), .ZN(n6460) );
NOR2_X1 U18913 ( .A1(n8677), .A2(n20882), .ZN(n8675) );
NOR2_X1 U18914 ( .A1(n8677), .A2(n20892), .ZN(n9539) );
NOR2_X1 U18915 ( .A1(n7657), .A2(n7658), .ZN(n7655) );
NOR2_X1 U18916 ( .A1(n8677), .A2(n20891), .ZN(n9252) );
NOR2_X1 U18917 ( .A1(n8677), .A2(n20887), .ZN(n9006) );
NOR2_X1 U18918 ( .A1(n20935), .A2(n6522), .ZN(n6520) );
NAND2_X1 U18919 ( .A1(n15797), .A2(n15916), .ZN(n6522) );
NOR2_X1 U18920 ( .A1(n7647), .A2(n20888), .ZN(n7645) );
NOR2_X1 U18921 ( .A1(n7649), .A2(n7650), .ZN(n7647) );
NAND2_X1 U18922 ( .A1(n7653), .A2(n7654), .ZN(n7649) );
OR2_X1 U18923 ( .A1(n7651), .A2(n20890), .ZN(n7650) );
NAND2_X1 U18924 ( .A1(n5898), .A2(n5899), .ZN(ex_block_i_alu_i_adder_in_b_31) );
NOR2_X1 U18925 ( .A1(n5912), .A2(n5913), .ZN(n5898) );
NOR2_X1 U18926 ( .A1(n5900), .A2(n5901), .ZN(n5899) );
NOR2_X1 U18927 ( .A1(n5917), .A2(n16095), .ZN(n5912) );
NAND2_X1 U18928 ( .A1(n6255), .A2(n6256), .ZN(ex_block_i_alu_i_adder_in_a_30) );
NAND2_X1 U18929 ( .A1(n6238), .A2(n15874), .ZN(n6255) );
NAND2_X1 U18930 ( .A1(n16357), .A2(n495), .ZN(n6256) );
NAND2_X1 U18931 ( .A1(n6253), .A2(n6254), .ZN(ex_block_i_alu_i_adder_in_a_31) );
NAND2_X1 U18932 ( .A1(n16408), .A2(n15875), .ZN(n6253) );
NAND2_X1 U18933 ( .A1(n16357), .A2(n414), .ZN(n6254) );
NAND2_X1 U18934 ( .A1(n9757), .A2(n9758), .ZN(n1275) );
NOR2_X1 U18935 ( .A1(n9774), .A2(n9775), .ZN(n9757) );
NOR2_X1 U18936 ( .A1(n9759), .A2(n9760), .ZN(n9758) );
NAND2_X1 U18937 ( .A1(n9785), .A2(n9786), .ZN(n9774) );
NAND2_X1 U18938 ( .A1(n9716), .A2(n9717), .ZN(n1236) );
NOR2_X1 U18939 ( .A1(n9730), .A2(n9731), .ZN(n9716) );
NOR2_X1 U18940 ( .A1(n9718), .A2(n9719), .ZN(n9717) );
NAND2_X1 U18941 ( .A1(n9732), .A2(n9733), .ZN(n9731) );
NAND2_X1 U18942 ( .A1(n9898), .A2(n9899), .ZN(n1415) );
NOR2_X1 U18943 ( .A1(n9930), .A2(n9931), .ZN(n9898) );
NOR2_X1 U18944 ( .A1(n9900), .A2(n9901), .ZN(n9899) );
NAND2_X1 U18945 ( .A1(n9939), .A2(n9940), .ZN(n9930) );
NAND2_X1 U18946 ( .A1(n9605), .A2(n9606), .ZN(n1119) );
NOR2_X1 U18947 ( .A1(n9618), .A2(n9619), .ZN(n9605) );
NOR2_X1 U18948 ( .A1(n9607), .A2(n9608), .ZN(n9606) );
NAND2_X1 U18949 ( .A1(n9620), .A2(n9621), .ZN(n9619) );
NAND2_X1 U18950 ( .A1(n9642), .A2(n9643), .ZN(n1158) );
NOR2_X1 U18951 ( .A1(n9655), .A2(n9656), .ZN(n9642) );
NOR2_X1 U18952 ( .A1(n9644), .A2(n9645), .ZN(n9643) );
NAND2_X1 U18953 ( .A1(n9657), .A2(n9658), .ZN(n9656) );
NAND2_X1 U18954 ( .A1(n9679), .A2(n9680), .ZN(n1197) );
NOR2_X1 U18955 ( .A1(n9692), .A2(n9693), .ZN(n9679) );
NOR2_X1 U18956 ( .A1(n9681), .A2(n9682), .ZN(n9680) );
NAND2_X1 U18957 ( .A1(n9694), .A2(n9695), .ZN(n9693) );
NAND2_X1 U18958 ( .A1(n9804), .A2(n9805), .ZN(n1331) );
NOR2_X1 U18959 ( .A1(n9817), .A2(n9818), .ZN(n9804) );
NOR2_X1 U18960 ( .A1(n9806), .A2(n9807), .ZN(n9805) );
NAND2_X1 U18961 ( .A1(n9819), .A2(n9820), .ZN(n9818) );
NAND2_X1 U18962 ( .A1(n6307), .A2(n6308), .ZN(ex_block_i_alu_i_shift_operand_31) );
NAND2_X1 U18963 ( .A1(n16467), .A2(n1391), .ZN(n6308) );
NAND2_X1 U18964 ( .A1(n1338), .A2(n5799), .ZN(n6307) );
NAND2_X1 U18965 ( .A1(n6517), .A2(n6518), .ZN(data_be_o_2_) );
NOR2_X1 U18966 ( .A1(n6523), .A2(n6524), .ZN(n6517) );
NOR2_X1 U18967 ( .A1(n6519), .A2(n6520), .ZN(n6518) );
NOR2_X1 U18968 ( .A1(n6526), .A2(n16407), .ZN(n6523) );
INV_X1 U18969 ( .A(n3442), .ZN(n20748) );
INV_X1 U18970 ( .A(n3427), .ZN(n20742) );
INV_X1 U18971 ( .A(n3422), .ZN(n20737) );
INV_X1 U18972 ( .A(n3417), .ZN(n20731) );
NAND2_X1 U18973 ( .A1(n6499), .A2(n6500), .ZN(data_wdata_o_0_) );
NOR2_X1 U18974 ( .A1(n6501), .A2(n6502), .ZN(n6500) );
NOR2_X1 U18975 ( .A1(n6503), .A2(n6504), .ZN(n6499) );
NOR2_X1 U18976 ( .A1(n20836), .A2(n16463), .ZN(n6501) );
NAND2_X1 U18977 ( .A1(n6433), .A2(n6434), .ZN(data_wdata_o_1_) );
NOR2_X1 U18978 ( .A1(n6435), .A2(n6436), .ZN(n6434) );
NOR2_X1 U18979 ( .A1(n6437), .A2(n6438), .ZN(n6433) );
NOR2_X1 U18980 ( .A1(n20834), .A2(n16463), .ZN(n6435) );
NAND2_X1 U18981 ( .A1(n6493), .A2(n6494), .ZN(data_wdata_o_10_) );
NOR2_X1 U18982 ( .A1(n6495), .A2(n6496), .ZN(n6494) );
NOR2_X1 U18983 ( .A1(n6497), .A2(n6498), .ZN(n6493) );
NOR2_X1 U18984 ( .A1(n20803), .A2(n16463), .ZN(n6495) );
NAND2_X1 U18985 ( .A1(n6487), .A2(n6488), .ZN(data_wdata_o_11_) );
NOR2_X1 U18986 ( .A1(n6489), .A2(n6490), .ZN(n6488) );
NOR2_X1 U18987 ( .A1(n6491), .A2(n6492), .ZN(n6487) );
NOR2_X1 U18988 ( .A1(n20800), .A2(n16463), .ZN(n6489) );
NAND2_X1 U18989 ( .A1(n6481), .A2(n6482), .ZN(data_wdata_o_12_) );
NOR2_X1 U18990 ( .A1(n6483), .A2(n6484), .ZN(n6482) );
NOR2_X1 U18991 ( .A1(n6485), .A2(n6486), .ZN(n6481) );
NOR2_X1 U18992 ( .A1(n20797), .A2(n16463), .ZN(n6483) );
NAND2_X1 U18993 ( .A1(n6475), .A2(n6476), .ZN(data_wdata_o_13_) );
NOR2_X1 U18994 ( .A1(n6477), .A2(n6478), .ZN(n6476) );
NOR2_X1 U18995 ( .A1(n6479), .A2(n6480), .ZN(n6475) );
NOR2_X1 U18996 ( .A1(n20794), .A2(n16463), .ZN(n6477) );
NAND2_X1 U18997 ( .A1(n6469), .A2(n6470), .ZN(data_wdata_o_14_) );
NOR2_X1 U18998 ( .A1(n6471), .A2(n6472), .ZN(n6470) );
NOR2_X1 U18999 ( .A1(n6473), .A2(n6474), .ZN(n6469) );
NOR2_X1 U19000 ( .A1(n20791), .A2(n16463), .ZN(n6471) );
NAND2_X1 U19001 ( .A1(n6463), .A2(n6464), .ZN(data_wdata_o_15_) );
NOR2_X1 U19002 ( .A1(n6465), .A2(n6466), .ZN(n6464) );
NOR2_X1 U19003 ( .A1(n6467), .A2(n6468), .ZN(n6463) );
NOR2_X1 U19004 ( .A1(n20788), .A2(n16463), .ZN(n6465) );
NAND2_X1 U19005 ( .A1(n6457), .A2(n6458), .ZN(data_wdata_o_16_) );
NOR2_X1 U19006 ( .A1(n6459), .A2(n6460), .ZN(n6458) );
NOR2_X1 U19007 ( .A1(n6461), .A2(n6462), .ZN(n6457) );
NOR2_X1 U19008 ( .A1(n20785), .A2(n16463), .ZN(n6459) );
NAND2_X1 U19009 ( .A1(n6451), .A2(n6452), .ZN(data_wdata_o_17_) );
NOR2_X1 U19010 ( .A1(n6453), .A2(n6454), .ZN(n6452) );
NOR2_X1 U19011 ( .A1(n6455), .A2(n6456), .ZN(n6451) );
NOR2_X1 U19012 ( .A1(n20782), .A2(n16463), .ZN(n6453) );
NAND2_X1 U19013 ( .A1(n6445), .A2(n6446), .ZN(data_wdata_o_18_) );
NOR2_X1 U19014 ( .A1(n6447), .A2(n6448), .ZN(n6446) );
NOR2_X1 U19015 ( .A1(n6449), .A2(n6450), .ZN(n6445) );
NOR2_X1 U19016 ( .A1(n20779), .A2(n16463), .ZN(n6447) );
NAND2_X1 U19017 ( .A1(n6439), .A2(n6440), .ZN(data_wdata_o_19_) );
NOR2_X1 U19018 ( .A1(n6441), .A2(n6442), .ZN(n6440) );
NOR2_X1 U19019 ( .A1(n6443), .A2(n6444), .ZN(n6439) );
NOR2_X1 U19020 ( .A1(n20776), .A2(n16463), .ZN(n6441) );
NAND2_X1 U19021 ( .A1(n6427), .A2(n6428), .ZN(data_wdata_o_20_) );
NOR2_X1 U19022 ( .A1(n6429), .A2(n6430), .ZN(n6428) );
NOR2_X1 U19023 ( .A1(n6431), .A2(n6432), .ZN(n6427) );
NOR2_X1 U19024 ( .A1(n20773), .A2(n16464), .ZN(n6429) );
NAND2_X1 U19025 ( .A1(n6421), .A2(n6422), .ZN(data_wdata_o_21_) );
NOR2_X1 U19026 ( .A1(n6423), .A2(n6424), .ZN(n6422) );
NOR2_X1 U19027 ( .A1(n6425), .A2(n6426), .ZN(n6421) );
NOR2_X1 U19028 ( .A1(n20770), .A2(n16464), .ZN(n6423) );
NAND2_X1 U19029 ( .A1(n6415), .A2(n6416), .ZN(data_wdata_o_22_) );
NOR2_X1 U19030 ( .A1(n6417), .A2(n6418), .ZN(n6416) );
NOR2_X1 U19031 ( .A1(n6419), .A2(n6420), .ZN(n6415) );
NOR2_X1 U19032 ( .A1(n20767), .A2(n16464), .ZN(n6417) );
NAND2_X1 U19033 ( .A1(n6409), .A2(n6410), .ZN(data_wdata_o_23_) );
NOR2_X1 U19034 ( .A1(n6411), .A2(n6412), .ZN(n6410) );
NOR2_X1 U19035 ( .A1(n6413), .A2(n6414), .ZN(n6409) );
NOR2_X1 U19036 ( .A1(n20764), .A2(n16464), .ZN(n6411) );
NAND2_X1 U19037 ( .A1(n6403), .A2(n6404), .ZN(data_wdata_o_24_) );
NOR2_X1 U19038 ( .A1(n6405), .A2(n6406), .ZN(n6404) );
NOR2_X1 U19039 ( .A1(n6407), .A2(n6408), .ZN(n6403) );
NOR2_X1 U19040 ( .A1(n20872), .A2(n16464), .ZN(n6405) );
NAND2_X1 U19041 ( .A1(n6397), .A2(n6398), .ZN(data_wdata_o_25_) );
NOR2_X1 U19042 ( .A1(n6399), .A2(n6400), .ZN(n6398) );
NOR2_X1 U19043 ( .A1(n6401), .A2(n6402), .ZN(n6397) );
NOR2_X1 U19044 ( .A1(n20870), .A2(n16464), .ZN(n6399) );
NAND2_X1 U19045 ( .A1(n6391), .A2(n6392), .ZN(data_wdata_o_26_) );
NOR2_X1 U19046 ( .A1(n6393), .A2(n6394), .ZN(n6392) );
NOR2_X1 U19047 ( .A1(n6395), .A2(n6396), .ZN(n6391) );
NOR2_X1 U19048 ( .A1(n20865), .A2(n16464), .ZN(n6393) );
NAND2_X1 U19049 ( .A1(n6385), .A2(n6386), .ZN(data_wdata_o_27_) );
NOR2_X1 U19050 ( .A1(n6387), .A2(n6388), .ZN(n6386) );
NOR2_X1 U19051 ( .A1(n6389), .A2(n6390), .ZN(n6385) );
NOR2_X1 U19052 ( .A1(n20862), .A2(n16464), .ZN(n6387) );
NAND2_X1 U19053 ( .A1(n6379), .A2(n6380), .ZN(data_wdata_o_28_) );
NOR2_X1 U19054 ( .A1(n6381), .A2(n6382), .ZN(n6380) );
NOR2_X1 U19055 ( .A1(n6383), .A2(n6384), .ZN(n6379) );
NOR2_X1 U19056 ( .A1(n20854), .A2(n16464), .ZN(n6381) );
NAND2_X1 U19057 ( .A1(n6373), .A2(n6374), .ZN(data_wdata_o_29_) );
NOR2_X1 U19058 ( .A1(n6375), .A2(n6376), .ZN(n6374) );
NOR2_X1 U19059 ( .A1(n6377), .A2(n6378), .ZN(n6373) );
NOR2_X1 U19060 ( .A1(n20847), .A2(n16464), .ZN(n6375) );
NOR2_X1 U19061 ( .A1(n10037), .A2(n10038), .ZN(n10030) );
NAND2_X1 U19062 ( .A1(n10039), .A2(n10040), .ZN(n10038) );
NAND2_X1 U19063 ( .A1(n10044), .A2(n10045), .ZN(n10037) );
NAND2_X1 U19064 ( .A1(alu_operand_b_ex_1), .A2(n10043), .ZN(n10039) );
NOR2_X1 U19065 ( .A1(n16254), .A2(n16255), .ZN(n16253) );
AND2_X1 U19066 ( .A1(n16468), .A2(n495), .ZN(n16254) );
AND2_X1 U19067 ( .A1(n16466), .A2(n466), .ZN(n16255) );
INV_X1 U19068 ( .A(n7603), .ZN(n20884) );
NAND2_X1 U19069 ( .A1(n9954), .A2(n9955), .ZN(n9782) );
NOR2_X1 U19070 ( .A1(n20838), .A2(n1297), .ZN(n9954) );
NOR2_X1 U19071 ( .A1(n20841), .A2(n20827), .ZN(n9955) );
NAND2_X1 U19072 ( .A1(alu_operand_b_ex_1), .A2(n20871), .ZN(n21649) );
AND2_X1 U19073 ( .A1(n7581), .A2(n7590), .ZN(n4020) );
NAND2_X1 U19074 ( .A1(n20884), .A2(n5128), .ZN(n7590) );
NAND2_X1 U19075 ( .A1(n9945), .A2(n20837), .ZN(n9924) );
NOR2_X1 U19076 ( .A1(n20827), .A2(n1297), .ZN(n9945) );
AND2_X1 U19077 ( .A1(n7581), .A2(n7671), .ZN(n3726) );
NAND2_X1 U19078 ( .A1(n7672), .A2(n20883), .ZN(n7671) );
NOR2_X1 U19079 ( .A1(n7619), .A2(n7685), .ZN(n7672) );
INV_X1 U19080 ( .A(n7656), .ZN(n20883) );
AND2_X1 U19081 ( .A1(n7581), .A2(n7598), .ZN(n4028) );
NAND2_X1 U19082 ( .A1(n7599), .A2(n20885), .ZN(n7598) );
NOR2_X1 U19083 ( .A1(n7601), .A2(n20893), .ZN(n7599) );
NOR2_X1 U19084 ( .A1(n7603), .A2(n7604), .ZN(n7601) );
NAND2_X1 U19085 ( .A1(n7674), .A2(n7675), .ZN(n7656) );
NOR2_X1 U19086 ( .A1(n7676), .A2(n7677), .ZN(n7674) );
NOR2_X1 U19087 ( .A1(n20893), .A2(n20884), .ZN(n7675) );
NOR2_X1 U19088 ( .A1(n20886), .A2(n7623), .ZN(n7677) );
NAND2_X1 U19089 ( .A1(n8896), .A2(n8897), .ZN(n383) );
NOR2_X1 U19090 ( .A1(n8898), .A2(n8899), .ZN(n8897) );
NOR2_X1 U19091 ( .A1(n8910), .A2(n8911), .ZN(n8896) );
NAND2_X1 U19092 ( .A1(n8900), .A2(n8901), .ZN(n8899) );
NAND2_X1 U19093 ( .A1(n8739), .A2(n8740), .ZN(n260) );
NOR2_X1 U19094 ( .A1(n8741), .A2(n8742), .ZN(n8740) );
NOR2_X1 U19095 ( .A1(n8754), .A2(n8755), .ZN(n8739) );
NAND2_X1 U19096 ( .A1(n8743), .A2(n8744), .ZN(n8742) );
NAND2_X1 U19097 ( .A1(n8701), .A2(n8702), .ZN(n218) );
NOR2_X1 U19098 ( .A1(n8714), .A2(n8715), .ZN(n8701) );
NOR2_X1 U19099 ( .A1(n8703), .A2(n8704), .ZN(n8702) );
NAND2_X1 U19100 ( .A1(n8716), .A2(n8717), .ZN(n8715) );
NAND2_X1 U19101 ( .A1(n9349), .A2(n9350), .ZN(n859) );
NOR2_X1 U19102 ( .A1(n9365), .A2(n9366), .ZN(n9349) );
NOR2_X1 U19103 ( .A1(n9351), .A2(n9352), .ZN(n9350) );
NAND2_X1 U19104 ( .A1(n9367), .A2(n9368), .ZN(n9366) );
NAND2_X1 U19105 ( .A1(n8932), .A2(n8933), .ZN(n427) );
NOR2_X1 U19106 ( .A1(n8948), .A2(n8949), .ZN(n8932) );
NOR2_X1 U19107 ( .A1(n8934), .A2(n8935), .ZN(n8933) );
NAND2_X1 U19108 ( .A1(n8950), .A2(n8951), .ZN(n8949) );
NAND2_X1 U19109 ( .A1(n9060), .A2(n9061), .ZN(n590) );
NOR2_X1 U19110 ( .A1(n9062), .A2(n9063), .ZN(n9061) );
NOR2_X1 U19111 ( .A1(n9076), .A2(n9077), .ZN(n9060) );
NAND2_X1 U19112 ( .A1(n9064), .A2(n9065), .ZN(n9063) );
NAND2_X1 U19113 ( .A1(n9101), .A2(n9102), .ZN(n630) );
NOR2_X1 U19114 ( .A1(n9103), .A2(n9104), .ZN(n9102) );
NOR2_X1 U19115 ( .A1(n9117), .A2(n9118), .ZN(n9101) );
NAND2_X1 U19116 ( .A1(n9105), .A2(n9106), .ZN(n9104) );
NAND2_X1 U19117 ( .A1(n9142), .A2(n9143), .ZN(n669) );
NOR2_X1 U19118 ( .A1(n9144), .A2(n9145), .ZN(n9143) );
NOR2_X1 U19119 ( .A1(n9158), .A2(n9159), .ZN(n9142) );
NAND2_X1 U19120 ( .A1(n9146), .A2(n9147), .ZN(n9145) );
NAND2_X1 U19121 ( .A1(n9183), .A2(n9184), .ZN(n707) );
NOR2_X1 U19122 ( .A1(n9185), .A2(n9186), .ZN(n9184) );
NOR2_X1 U19123 ( .A1(n9199), .A2(n9200), .ZN(n9183) );
NAND2_X1 U19124 ( .A1(n9187), .A2(n9188), .ZN(n9186) );
NAND2_X1 U19125 ( .A1(n9224), .A2(n9225), .ZN(n744) );
NOR2_X1 U19126 ( .A1(n9226), .A2(n9227), .ZN(n9225) );
NOR2_X1 U19127 ( .A1(n9240), .A2(n9241), .ZN(n9224) );
NAND2_X1 U19128 ( .A1(n9228), .A2(n9229), .ZN(n9227) );
NAND2_X1 U19129 ( .A1(n9265), .A2(n9266), .ZN(n782) );
NOR2_X1 U19130 ( .A1(n9267), .A2(n9268), .ZN(n9266) );
NOR2_X1 U19131 ( .A1(n9281), .A2(n9282), .ZN(n9265) );
NAND2_X1 U19132 ( .A1(n9269), .A2(n9270), .ZN(n9268) );
NAND2_X1 U19133 ( .A1(n9436), .A2(n9437), .ZN(n940) );
NOR2_X1 U19134 ( .A1(n9438), .A2(n9439), .ZN(n9437) );
NOR2_X1 U19135 ( .A1(n9452), .A2(n9453), .ZN(n9436) );
NAND2_X1 U19136 ( .A1(n9440), .A2(n9441), .ZN(n9439) );
NAND2_X1 U19137 ( .A1(n9477), .A2(n9478), .ZN(n979) );
NOR2_X1 U19138 ( .A1(n9479), .A2(n9480), .ZN(n9478) );
NOR2_X1 U19139 ( .A1(n9493), .A2(n9494), .ZN(n9477) );
NAND2_X1 U19140 ( .A1(n9481), .A2(n9482), .ZN(n9480) );
NAND2_X1 U19141 ( .A1(n9563), .A2(n9564), .ZN(n1075) );
NOR2_X1 U19142 ( .A1(n9565), .A2(n9566), .ZN(n9564) );
NOR2_X1 U19143 ( .A1(n9579), .A2(n9580), .ZN(n9563) );
NAND2_X1 U19144 ( .A1(n9567), .A2(n9568), .ZN(n9566) );
NAND2_X1 U19145 ( .A1(n8558), .A2(n8559), .ZN(n79) );
NOR2_X1 U19146 ( .A1(n8577), .A2(n8578), .ZN(n8558) );
NOR2_X1 U19147 ( .A1(n8560), .A2(n8561), .ZN(n8559) );
NAND2_X1 U19148 ( .A1(n8579), .A2(n8580), .ZN(n8578) );
NAND2_X1 U19149 ( .A1(n8610), .A2(n8611), .ZN(n127) );
NOR2_X1 U19150 ( .A1(n8625), .A2(n8626), .ZN(n8610) );
NOR2_X1 U19151 ( .A1(n8612), .A2(n8613), .ZN(n8611) );
NAND2_X1 U19152 ( .A1(n8627), .A2(n8628), .ZN(n8626) );
NAND2_X1 U19153 ( .A1(n8783), .A2(n8784), .ZN(n301) );
NOR2_X1 U19154 ( .A1(n8785), .A2(n8786), .ZN(n8784) );
NOR2_X1 U19155 ( .A1(n8799), .A2(n8800), .ZN(n8783) );
NAND2_X1 U19156 ( .A1(n8787), .A2(n8788), .ZN(n8786) );
NAND2_X1 U19157 ( .A1(n8653), .A2(n8654), .ZN(n175) );
NOR2_X1 U19158 ( .A1(n8671), .A2(n8672), .ZN(n8653) );
NOR2_X1 U19159 ( .A1(n8655), .A2(n8656), .ZN(n8654) );
NAND2_X1 U19160 ( .A1(n8681), .A2(n8682), .ZN(n8671) );
NAND2_X1 U19161 ( .A1(n9852), .A2(n9853), .ZN(n472) );
NOR2_X1 U19162 ( .A1(n9871), .A2(n9872), .ZN(n9852) );
NOR2_X1 U19163 ( .A1(n9854), .A2(n9855), .ZN(n9853) );
NAND2_X1 U19164 ( .A1(n9879), .A2(n9880), .ZN(n9871) );
NAND2_X1 U19165 ( .A1(n9392), .A2(n9393), .ZN(n904) );
NOR2_X1 U19166 ( .A1(n9408), .A2(n9409), .ZN(n9392) );
NOR2_X1 U19167 ( .A1(n9394), .A2(n9395), .ZN(n9393) );
NAND2_X1 U19168 ( .A1(n9416), .A2(n9417), .ZN(n9408) );
NAND2_X1 U19169 ( .A1(n9019), .A2(n9020), .ZN(n550) );
NOR2_X1 U19170 ( .A1(n9021), .A2(n9022), .ZN(n9020) );
NOR2_X1 U19171 ( .A1(n9035), .A2(n9036), .ZN(n9019) );
NAND2_X1 U19172 ( .A1(n9023), .A2(n9024), .ZN(n9022) );
NAND2_X1 U19173 ( .A1(n8978), .A2(n8979), .ZN(n510) );
NOR2_X1 U19174 ( .A1(n8980), .A2(n8981), .ZN(n8979) );
NOR2_X1 U19175 ( .A1(n8994), .A2(n8995), .ZN(n8978) );
NAND2_X1 U19176 ( .A1(n8982), .A2(n8983), .ZN(n8981) );
NAND2_X1 U19177 ( .A1(n9306), .A2(n9307), .ZN(n820) );
NOR2_X1 U19178 ( .A1(n9323), .A2(n9324), .ZN(n9306) );
NOR2_X1 U19179 ( .A1(n9308), .A2(n9309), .ZN(n9307) );
NAND2_X1 U19180 ( .A1(n9331), .A2(n9332), .ZN(n9323) );
NAND2_X1 U19181 ( .A1(n9518), .A2(n9519), .ZN(n1017) );
NOR2_X1 U19182 ( .A1(n9535), .A2(n9536), .ZN(n9518) );
NOR2_X1 U19183 ( .A1(n9520), .A2(n9521), .ZN(n9519) );
NAND2_X1 U19184 ( .A1(n9544), .A2(n9545), .ZN(n9535) );
NAND2_X1 U19185 ( .A1(n8829), .A2(n8830), .ZN(n342) );
NOR2_X1 U19186 ( .A1(n8848), .A2(n8849), .ZN(n8829) );
NOR2_X1 U19187 ( .A1(n8831), .A2(n8832), .ZN(n8830) );
NAND2_X1 U19188 ( .A1(n8850), .A2(n8851), .ZN(n8849) );
NAND2_X1 U19189 ( .A1(n5918), .A2(n5919), .ZN(ex_block_i_alu_i_adder_in_b_30) );
NOR2_X1 U19190 ( .A1(n5928), .A2(n5929), .ZN(n5918) );
NOR2_X1 U19191 ( .A1(n5920), .A2(n5921), .ZN(n5919) );
NOR2_X1 U19192 ( .A1(n5917), .A2(n16096), .ZN(n5928) );
NAND2_X1 U19193 ( .A1(alu_operand_b_ex_2), .A2(n10002), .ZN(n10035) );
OR2_X1 U19194 ( .A1(alu_operand_b_ex_1), .A2(ex_block_i_alu_i_shift_amt_compl_0), .ZN(n21653) );
NAND2_X1 U19195 ( .A1(n8667), .A2(n16361), .ZN(n8666) );
NAND2_X1 U19196 ( .A1(n16386), .A2(n15974), .ZN(n8667) );
NAND2_X1 U19197 ( .A1(n20838), .A2(alu_operand_b_ex_3), .ZN(n9997) );
NAND2_X1 U19198 ( .A1(n10123), .A2(n10124), .ZN(n10116) );
OR2_X1 U19199 ( .A1(n5799), .A2(n10125), .ZN(n10124) );
NAND2_X1 U19200 ( .A1(n10125), .A2(n5799), .ZN(n10123) );
NOR2_X1 U19201 ( .A1(n20941), .A2(n10117), .ZN(n10125) );
NAND2_X1 U19202 ( .A1(n21658), .A2(n21657), .ZN(n21659) );
NOR2_X1 U19203 ( .A1(alu_operand_b_ex_1), .A2(ex_block_i_alu_i_shift_amt_compl_0), .ZN(n21658) );
NOR2_X1 U19204 ( .A1(alu_operand_b_ex_3), .A2(alu_operand_b_ex_2), .ZN(n21657) );
NAND2_X1 U19205 ( .A1(n16468), .A2(n5799), .ZN(n5797) );
NAND2_X1 U19206 ( .A1(n1338), .A2(n615), .ZN(n5761) );
NAND2_X1 U19207 ( .A1(n16467), .A2(n240), .ZN(n5762) );
NAND2_X1 U19208 ( .A1(n16466), .A2(n575), .ZN(n5759) );
NAND2_X1 U19209 ( .A1(n16468), .A2(n282), .ZN(n5760) );
NAND2_X1 U19210 ( .A1(n1338), .A2(n535), .ZN(n5757) );
NAND2_X1 U19211 ( .A1(n16468), .A2(n323), .ZN(n5758) );
NAND2_X1 U19212 ( .A1(n16468), .A2(n51), .ZN(n5769) );
NAND2_X1 U19213 ( .A1(n1338), .A2(n768), .ZN(n5770) );
NAND2_X1 U19214 ( .A1(n16468), .A2(n883), .ZN(n5751) );
NAND2_X1 U19215 ( .A1(n1338), .A2(n414), .ZN(n5752) );
NAND2_X1 U19216 ( .A1(n16466), .A2(n845), .ZN(n5774) );
NAND2_X1 U19217 ( .A1(n16467), .A2(n1258), .ZN(n5773) );
NAND2_X1 U19218 ( .A1(n16467), .A2(n535), .ZN(n5749) );
NAND2_X1 U19219 ( .A1(n1338), .A2(n323), .ZN(n5750) );
NAND2_X1 U19220 ( .A1(n16468), .A2(n575), .ZN(n5747) );
NAND2_X1 U19221 ( .A1(n16466), .A2(n282), .ZN(n5748) );
NAND2_X1 U19222 ( .A1(n16467), .A2(n615), .ZN(n5745) );
NAND2_X1 U19223 ( .A1(n1338), .A2(n240), .ZN(n5746) );
NAND2_X1 U19224 ( .A1(n16468), .A2(n655), .ZN(n5743) );
NAND2_X1 U19225 ( .A1(n16466), .A2(n213), .ZN(n5744) );
NAND2_X1 U19226 ( .A1(n16467), .A2(n1178), .ZN(n5779) );
NAND2_X1 U19227 ( .A1(n16466), .A2(n965), .ZN(n5780) );
NAND2_X1 U19228 ( .A1(n16467), .A2(n1139), .ZN(n5781) );
NAND2_X1 U19229 ( .A1(n1338), .A2(n1003), .ZN(n5782) );
INV_X1 U19230 ( .A(n412), .ZN(n20766) );
NAND2_X1 U19231 ( .A1(n7684), .A2(n7683), .ZN(n10343) );
NOR2_X1 U19232 ( .A1(n16257), .A2(n16258), .ZN(n16256) );
AND2_X1 U19233 ( .A1(n16466), .A2(n883), .ZN(n16257) );
AND2_X1 U19234 ( .A1(n16468), .A2(n414), .ZN(n16258) );
NAND2_X1 U19235 ( .A1(n1338), .A2(n495), .ZN(n5755) );
NAND2_X1 U19236 ( .A1(n16467), .A2(n466), .ZN(n5756) );
NAND2_X1 U19237 ( .A1(n1338), .A2(n655), .ZN(n5763) );
NAND2_X1 U19238 ( .A1(n16467), .A2(n213), .ZN(n5764) );
NAND2_X1 U19239 ( .A1(n1338), .A2(n693), .ZN(n5765) );
NAND2_X1 U19240 ( .A1(n16468), .A2(n170), .ZN(n5766) );
NAND2_X1 U19241 ( .A1(n16466), .A2(n730), .ZN(n5767) );
NAND2_X1 U19242 ( .A1(n16467), .A2(n107), .ZN(n5768) );
NAND2_X1 U19243 ( .A1(n1338), .A2(n1217), .ZN(n5791) );
NAND2_X1 U19244 ( .A1(n16468), .A2(n926), .ZN(n5792) );
NAND2_X1 U19245 ( .A1(n1338), .A2(n1102), .ZN(n5785) );
NAND2_X1 U19246 ( .A1(n16468), .A2(n1046), .ZN(n5786) );
NAND2_X1 U19247 ( .A1(n16466), .A2(n1139), .ZN(n5787) );
NAND2_X1 U19248 ( .A1(n16468), .A2(n1003), .ZN(n5788) );
NAND2_X1 U19249 ( .A1(n1338), .A2(n1178), .ZN(n5789) );
NAND2_X1 U19250 ( .A1(n16468), .A2(n965), .ZN(n5790) );
NAND2_X1 U19251 ( .A1(n15802), .A2(n15858), .ZN(n6514) );
NAND2_X1 U19252 ( .A1(n16466), .A2(n51), .ZN(n5737) );
NAND2_X1 U19253 ( .A1(n16467), .A2(n768), .ZN(n5738) );
NAND2_X1 U19254 ( .A1(n10025), .A2(n10026), .ZN(n10017) );
NAND2_X1 U19255 ( .A1(n20845), .A2(n20827), .ZN(n10025) );
NAND2_X1 U19256 ( .A1(n10027), .A2(n1297), .ZN(n10026) );
NAND2_X1 U19257 ( .A1(n10030), .A2(n10031), .ZN(n10027) );
NAND2_X1 U19258 ( .A1(n16467), .A2(n845), .ZN(n5794) );
NAND2_X1 U19259 ( .A1(n1338), .A2(n1258), .ZN(n5793) );
NAND2_X1 U19260 ( .A1(n1338), .A2(n1295), .ZN(n5795) );
NAND2_X1 U19261 ( .A1(n16467), .A2(n806), .ZN(n5796) );
OR2_X1 U19262 ( .A1(n21653), .A2(alu_operand_b_ex_2), .ZN(n21654) );
NAND2_X1 U19263 ( .A1(n5922), .A2(n5923), .ZN(n5921) );
NAND2_X1 U19264 ( .A1(n497), .A2(n5904), .ZN(n5922) );
NAND2_X1 U19265 ( .A1(n20769), .A2(n16409), .ZN(n5923) );
INV_X1 U19266 ( .A(n497), .ZN(n20769) );
NAND2_X1 U19267 ( .A1(n5902), .A2(n5903), .ZN(n5901) );
NAND2_X1 U19268 ( .A1(n412), .A2(n16334), .ZN(n5902) );
NAND2_X1 U19269 ( .A1(n20766), .A2(n5826), .ZN(n5903) );
NAND2_X1 U19270 ( .A1(ex_block_i_alu_i_adder_in_b_1), .A2(n16334), .ZN(n21131) );
NAND2_X1 U19271 ( .A1(n7626), .A2(n7627), .ZN(n7625) );
NAND2_X1 U19272 ( .A1(n20885), .A2(n7629), .ZN(n7626) );
NAND2_X1 U19273 ( .A1(n7628), .A2(n20884), .ZN(n7627) );
NAND2_X1 U19274 ( .A1(n9767), .A2(n9768), .ZN(n9759) );
NOR2_X1 U19275 ( .A1(n9769), .A2(n9770), .ZN(n9768) );
NOR2_X1 U19276 ( .A1(n9772), .A2(n9773), .ZN(n9767) );
NAND2_X1 U19277 ( .A1(n9771), .A2(n16361), .ZN(n9770) );
NAND2_X1 U19278 ( .A1(n9316), .A2(n9317), .ZN(n9308) );
NOR2_X1 U19279 ( .A1(n9318), .A2(n9319), .ZN(n9317) );
NOR2_X1 U19280 ( .A1(n9321), .A2(n9322), .ZN(n9316) );
NAND2_X1 U19281 ( .A1(n9320), .A2(n16361), .ZN(n9319) );
NAND2_X1 U19282 ( .A1(n9528), .A2(n9529), .ZN(n9520) );
NOR2_X1 U19283 ( .A1(n9530), .A2(n9531), .ZN(n9529) );
NOR2_X1 U19284 ( .A1(n9533), .A2(n9534), .ZN(n9528) );
NAND2_X1 U19285 ( .A1(n9532), .A2(n16361), .ZN(n9531) );
NAND2_X1 U19286 ( .A1(n7641), .A2(n7642), .ZN(n7640) );
NOR2_X1 U19287 ( .A1(n7643), .A2(n7644), .ZN(n7642) );
NOR2_X1 U19288 ( .A1(n7655), .A2(n7656), .ZN(n7641) );
NOR2_X1 U19289 ( .A1(n7645), .A2(n7646), .ZN(n7644) );
NAND2_X1 U19290 ( .A1(ex_block_i_alu_i_adder_in_b_2), .A2(n20754), .ZN(n21226) );
NAND2_X1 U19291 ( .A1(ex_block_i_alu_i_adder_in_b_3), .A2(n20750), .ZN(n21260) );
NAND2_X1 U19292 ( .A1(ex_block_i_alu_i_adder_in_b_4), .A2(n20744), .ZN(n21266) );
NAND2_X1 U19293 ( .A1(ex_block_i_alu_i_adder_in_b_5), .A2(n20739), .ZN(n21272) );
NAND2_X1 U19294 ( .A1(ex_block_i_alu_i_adder_in_b_6), .A2(n20733), .ZN(n21278) );
NAND2_X1 U19295 ( .A1(ex_block_i_alu_i_adder_in_b_7), .A2(n20728), .ZN(n21284) );
NAND2_X1 U19296 ( .A1(ex_block_i_alu_i_adder_in_b_8), .A2(n20722), .ZN(n21290) );
NAND2_X1 U19297 ( .A1(ex_block_i_alu_i_adder_in_b_9), .A2(n20717), .ZN(n21296) );
NAND2_X1 U19298 ( .A1(ex_block_i_alu_i_adder_in_b_10), .A2(n20713), .ZN(n21045) );
NAND2_X1 U19299 ( .A1(ex_block_i_alu_i_adder_in_b_11), .A2(n20709), .ZN(n21054) );
NAND2_X1 U19300 ( .A1(ex_block_i_alu_i_adder_in_b_12), .A2(n20705), .ZN(n21063) );
AND2_X1 U19301 ( .A1(n21653), .A2(alu_operand_b_ex_2), .ZN(n21652) );
AND2_X1 U19302 ( .A1(n21654), .A2(alu_operand_b_ex_3), .ZN(n21656) );
AND2_X1 U19303 ( .A1(n21659), .A2(alu_operand_b_ex_4), .ZN(n21661) );
NAND2_X1 U19304 ( .A1(ex_block_i_alu_i_adder_in_b_32), .A2(n16259), .ZN(n21250) );
AND2_X1 U19305 ( .A1(n9949), .A2(n9950), .ZN(n8581) );
NOR2_X1 U19306 ( .A1(n20845), .A2(n9952), .ZN(n9950) );
NOR2_X1 U19307 ( .A1(n7311), .A2(n9953), .ZN(n9949) );
NAND2_X1 U19308 ( .A1(n1297), .A2(alu_operand_b_ex_4), .ZN(n9952) );
NAND2_X1 U19309 ( .A1(n16386), .A2(n15976), .ZN(n9771) );
NAND2_X1 U19310 ( .A1(n16386), .A2(n15973), .ZN(n9320) );
NAND2_X1 U19311 ( .A1(n16386), .A2(n15975), .ZN(n9532) );
NOR2_X1 U19312 ( .A1(n16260), .A2(n16261), .ZN(n16259) );
AND2_X1 U19313 ( .A1(n20961), .A2(n5799), .ZN(n16260) );
AND2_X1 U19314 ( .A1(n16408), .A2(n15891), .ZN(n16261) );
OR2_X1 U19315 ( .A1(n20871), .A2(alu_operand_b_ex_1), .ZN(n21650) );
OR2_X1 U19316 ( .A1(n8121), .A2(n197), .ZN(n10040) );
OR2_X1 U19317 ( .A1(n5904), .A2(ex_block_i_alu_i_adder_in_b_1), .ZN(n21132) );
OR2_X1 U19318 ( .A1(n20744), .A2(ex_block_i_alu_i_adder_in_b_4), .ZN(n21267) );
OR2_X1 U19319 ( .A1(n20728), .A2(ex_block_i_alu_i_adder_in_b_7), .ZN(n21285) );
OR2_X1 U19320 ( .A1(n20722), .A2(ex_block_i_alu_i_adder_in_b_8), .ZN(n21291) );
OR2_X1 U19321 ( .A1(n20709), .A2(ex_block_i_alu_i_adder_in_b_11), .ZN(n21055) );
OR2_X1 U19322 ( .A1(n20754), .A2(ex_block_i_alu_i_adder_in_b_2), .ZN(n21227) );
OR2_X1 U19323 ( .A1(n20750), .A2(ex_block_i_alu_i_adder_in_b_3), .ZN(n21261) );
OR2_X1 U19324 ( .A1(n20739), .A2(ex_block_i_alu_i_adder_in_b_5), .ZN(n21273) );
OR2_X1 U19325 ( .A1(n20733), .A2(ex_block_i_alu_i_adder_in_b_6), .ZN(n21279) );
OR2_X1 U19326 ( .A1(n20717), .A2(ex_block_i_alu_i_adder_in_b_9), .ZN(n21297) );
OR2_X1 U19327 ( .A1(n20713), .A2(ex_block_i_alu_i_adder_in_b_10), .ZN(n21046) );
OR2_X1 U19328 ( .A1(n20705), .A2(ex_block_i_alu_i_adder_in_b_12), .ZN(n21064) );
OR2_X1 U19329 ( .A1(n16259), .A2(ex_block_i_alu_i_adder_in_b_32), .ZN(n21251) );
NAND2_X1 U19330 ( .A1(n1757), .A2(n1758), .ZN(instr_addr_o_2_) );
NAND2_X1 U19331 ( .A1(n15929), .A2(n15934), .ZN(n1758) );
NOR2_X1 U19332 ( .A1(n1760), .A2(n1761), .ZN(n1757) );
NOR2_X1 U19333 ( .A1(n20748), .A2(n1708), .ZN(n1760) );
NAND2_X1 U19334 ( .A1(n1739), .A2(n1740), .ZN(instr_addr_o_3_) );
NAND2_X1 U19335 ( .A1(n15929), .A2(n15935), .ZN(n1740) );
NOR2_X1 U19336 ( .A1(n1742), .A2(n1743), .ZN(n1739) );
NOR2_X1 U19337 ( .A1(n20742), .A2(n1708), .ZN(n1742) );
NAND2_X1 U19338 ( .A1(n1733), .A2(n1734), .ZN(instr_addr_o_4_) );
NAND2_X1 U19339 ( .A1(n15929), .A2(n15936), .ZN(n1734) );
NOR2_X1 U19340 ( .A1(n1736), .A2(n1737), .ZN(n1733) );
NOR2_X1 U19341 ( .A1(n20737), .A2(n1708), .ZN(n1736) );
NAND2_X1 U19342 ( .A1(n6527), .A2(n6528), .ZN(data_be_o_1_) );
OR2_X1 U19343 ( .A1(n6525), .A2(n1566), .ZN(n6528) );
NOR2_X1 U19344 ( .A1(n6529), .A2(n6530), .ZN(n6527) );
NOR2_X1 U19345 ( .A1(n6526), .A2(n16405), .ZN(n6530) );
NAND2_X1 U19346 ( .A1(n6367), .A2(n6368), .ZN(data_wdata_o_2_) );
NOR2_X1 U19347 ( .A1(n6369), .A2(n6370), .ZN(n6368) );
NOR2_X1 U19348 ( .A1(n6371), .A2(n6372), .ZN(n6367) );
NOR2_X1 U19349 ( .A1(n20831), .A2(n16464), .ZN(n6369) );
NAND2_X1 U19350 ( .A1(n6349), .A2(n6350), .ZN(data_wdata_o_3_) );
NOR2_X1 U19351 ( .A1(n6351), .A2(n6352), .ZN(n6350) );
NOR2_X1 U19352 ( .A1(n6353), .A2(n6354), .ZN(n6349) );
NOR2_X1 U19353 ( .A1(n20829), .A2(n16463), .ZN(n6351) );
NAND2_X1 U19354 ( .A1(n6343), .A2(n6344), .ZN(data_wdata_o_4_) );
NOR2_X1 U19355 ( .A1(n6345), .A2(n6346), .ZN(n6344) );
NOR2_X1 U19356 ( .A1(n6347), .A2(n6348), .ZN(n6343) );
NOR2_X1 U19357 ( .A1(n20817), .A2(n16464), .ZN(n6345) );
NAND2_X1 U19358 ( .A1(n6337), .A2(n6338), .ZN(data_wdata_o_5_) );
NOR2_X1 U19359 ( .A1(n6339), .A2(n6340), .ZN(n6338) );
NOR2_X1 U19360 ( .A1(n6341), .A2(n6342), .ZN(n6337) );
NOR2_X1 U19361 ( .A1(n20815), .A2(n16463), .ZN(n6339) );
NAND2_X1 U19362 ( .A1(n6331), .A2(n6332), .ZN(data_wdata_o_6_) );
NOR2_X1 U19363 ( .A1(n6333), .A2(n6334), .ZN(n6332) );
NOR2_X1 U19364 ( .A1(n6335), .A2(n6336), .ZN(n6331) );
NOR2_X1 U19365 ( .A1(n20813), .A2(n16464), .ZN(n6333) );
NAND2_X1 U19366 ( .A1(n6325), .A2(n6326), .ZN(data_wdata_o_7_) );
NOR2_X1 U19367 ( .A1(n6327), .A2(n6328), .ZN(n6326) );
NOR2_X1 U19368 ( .A1(n6329), .A2(n6330), .ZN(n6325) );
NOR2_X1 U19369 ( .A1(n20811), .A2(n16463), .ZN(n6327) );
NAND2_X1 U19370 ( .A1(n6319), .A2(n6320), .ZN(data_wdata_o_8_) );
NOR2_X1 U19371 ( .A1(n6321), .A2(n6322), .ZN(n6320) );
NOR2_X1 U19372 ( .A1(n6323), .A2(n6324), .ZN(n6319) );
NOR2_X1 U19373 ( .A1(n20809), .A2(n16464), .ZN(n6321) );
NAND2_X1 U19374 ( .A1(n6311), .A2(n6312), .ZN(data_wdata_o_9_) );
NOR2_X1 U19375 ( .A1(n6313), .A2(n6314), .ZN(n6312) );
NOR2_X1 U19376 ( .A1(n6316), .A2(n6317), .ZN(n6311) );
NOR2_X1 U19377 ( .A1(n20806), .A2(n16463), .ZN(n6313) );
NAND2_X1 U19378 ( .A1(n6361), .A2(n6362), .ZN(data_wdata_o_30_) );
NOR2_X1 U19379 ( .A1(n6363), .A2(n6364), .ZN(n6362) );
NOR2_X1 U19380 ( .A1(n6365), .A2(n6366), .ZN(n6361) );
NOR2_X1 U19381 ( .A1(n20842), .A2(n16464), .ZN(n6363) );
NAND2_X1 U19382 ( .A1(n6355), .A2(n6356), .ZN(data_wdata_o_31_) );
NOR2_X1 U19383 ( .A1(n6357), .A2(n6358), .ZN(n6356) );
NOR2_X1 U19384 ( .A1(n6359), .A2(n6360), .ZN(n6355) );
NOR2_X1 U19385 ( .A1(n20840), .A2(n16464), .ZN(n6357) );
NAND2_X1 U19386 ( .A1(n6533), .A2(n6534), .ZN(data_be_o_0_) );
NOR2_X1 U19387 ( .A1(n6519), .A2(n6529), .ZN(n6534) );
NOR2_X1 U19388 ( .A1(n6538), .A2(n6539), .ZN(n6533) );
NOR2_X1 U19389 ( .A1(n6540), .A2(n1566), .ZN(n6539) );
NAND2_X1 U19390 ( .A1(n1038), .A2(n1039), .ZN(n376) );
NOR2_X1 U19391 ( .A1(n1040), .A2(n33), .ZN(n1038) );
NAND2_X1 U19392 ( .A1(n1365), .A2(n1366), .ZN(n33) );
NOR2_X1 U19393 ( .A1(n19989), .A2(n1368), .ZN(n1366) );
NAND2_X1 U19394 ( .A1(n20993), .A2(n20022), .ZN(n1368) );
NOR2_X1 U19395 ( .A1(n20000), .A2(n378), .ZN(n499) );
NOR2_X1 U19396 ( .A1(n19999), .A2(n378), .ZN(n416) );
NOR2_X1 U19397 ( .A1(n373), .A2(n374), .ZN(n365) );
NOR2_X1 U19398 ( .A1(n19998), .A2(n378), .ZN(n373) );
NOR2_X1 U19399 ( .A1(n19990), .A2(n376), .ZN(n374) );
NOR2_X1 U19400 ( .A1(n65), .A2(n16335), .ZN(n55) );
NOR2_X1 U19401 ( .A1(n66), .A2(n67), .ZN(n65) );
NAND2_X1 U19402 ( .A1(n68), .A2(n69), .ZN(n67) );
NOR2_X1 U19403 ( .A1(n72), .A2(n20004), .ZN(n66) );
NOR2_X1 U19404 ( .A1(n117), .A2(n33), .ZN(n110) );
NOR2_X1 U19405 ( .A1(n118), .A2(n119), .ZN(n117) );
NAND2_X1 U19406 ( .A1(n120), .A2(n121), .ZN(n119) );
NOR2_X1 U19407 ( .A1(n72), .A2(n20005), .ZN(n118) );
NOR2_X1 U19408 ( .A1(n890), .A2(n16335), .ZN(n889) );
NOR2_X1 U19409 ( .A1(n891), .A2(n892), .ZN(n890) );
NAND2_X1 U19410 ( .A1(n895), .A2(n896), .ZN(n891) );
NAND2_X1 U19411 ( .A1(n893), .A2(n894), .ZN(n892) );
NOR2_X1 U19412 ( .A1(n330), .A2(n16335), .ZN(n329) );
NOR2_X1 U19413 ( .A1(n331), .A2(n332), .ZN(n330) );
NAND2_X1 U19414 ( .A1(n335), .A2(n336), .ZN(n331) );
NAND2_X1 U19415 ( .A1(n333), .A2(n334), .ZN(n332) );
NOR2_X1 U19416 ( .A1(n289), .A2(n33), .ZN(n288) );
NOR2_X1 U19417 ( .A1(n290), .A2(n291), .ZN(n289) );
NAND2_X1 U19418 ( .A1(n294), .A2(n295), .ZN(n290) );
NAND2_X1 U19419 ( .A1(n292), .A2(n293), .ZN(n291) );
NOR2_X1 U19420 ( .A1(n20006), .A2(n44), .ZN(n360) );
NOR2_X1 U19421 ( .A1(n725), .A2(n726), .ZN(n722) );
NOR2_X1 U19422 ( .A1(n19998), .A2(n376), .ZN(n725) );
NOR2_X1 U19423 ( .A1(n20014), .A2(n16477), .ZN(n726) );
INV_X1 U19424 ( .A(n1391), .ZN(n20759) );
NOR2_X1 U19425 ( .A1(n1058), .A2(n19990), .ZN(n1306) );
NOR2_X1 U19426 ( .A1(n7620), .A2(n7621), .ZN(n7617) );
NAND2_X1 U19427 ( .A1(n7622), .A2(n7623), .ZN(n7621) );
NOR2_X1 U19428 ( .A1(n20005), .A2(n897), .ZN(n1357) );
NOR2_X1 U19429 ( .A1(n1040), .A2(n20014), .ZN(n1307) );
NOR2_X1 U19430 ( .A1(n1040), .A2(n20021), .ZN(n1363) );
NOR2_X1 U19431 ( .A1(n20013), .A2(n898), .ZN(n1358) );
INV_X1 U19432 ( .A(n466), .ZN(n20751) );
INV_X1 U19433 ( .A(n213), .ZN(n20729) );
INV_X1 U19434 ( .A(n170), .ZN(n20723) );
NOR2_X1 U19435 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NOR2_X1 U19436 ( .A1(n1304), .A2(n20006), .ZN(n1303) );
NOR2_X1 U19437 ( .A1(n1305), .A2(n19998), .ZN(n1302) );
NOR2_X1 U19438 ( .A1(n1036), .A2(n1037), .ZN(n1033) );
NOR2_X1 U19439 ( .A1(n44), .A2(n20021), .ZN(n1037) );
NOR2_X1 U19440 ( .A1(n20005), .A2(n376), .ZN(n1036) );
NOR2_X1 U19441 ( .A1(n998), .A2(n999), .ZN(n995) );
NOR2_X1 U19442 ( .A1(n20004), .A2(n376), .ZN(n998) );
NOR2_X1 U19443 ( .A1(n20020), .A2(n16477), .ZN(n999) );
NOR2_X1 U19444 ( .A1(n920), .A2(n921), .ZN(n917) );
NOR2_X1 U19445 ( .A1(n44), .A2(n20018), .ZN(n921) );
NOR2_X1 U19446 ( .A1(n20002), .A2(n376), .ZN(n920) );
NOR2_X1 U19447 ( .A1(n839), .A2(n840), .ZN(n836) );
NOR2_X1 U19448 ( .A1(n44), .A2(n20017), .ZN(n840) );
NOR2_X1 U19449 ( .A1(n20001), .A2(n376), .ZN(n839) );
NOR2_X1 U19450 ( .A1(n800), .A2(n801), .ZN(n797) );
NOR2_X1 U19451 ( .A1(n44), .A2(n20016), .ZN(n801) );
NOR2_X1 U19452 ( .A1(n20000), .A2(n376), .ZN(n800) );
NOR2_X1 U19453 ( .A1(n762), .A2(n763), .ZN(n759) );
NOR2_X1 U19454 ( .A1(n44), .A2(n20015), .ZN(n763) );
NOR2_X1 U19455 ( .A1(n19999), .A2(n376), .ZN(n762) );
NOR2_X1 U19456 ( .A1(n959), .A2(n960), .ZN(n956) );
NOR2_X1 U19457 ( .A1(n44), .A2(n20019), .ZN(n960) );
NOR2_X1 U19458 ( .A1(n376), .A2(n20003), .ZN(n959) );
NAND2_X1 U19459 ( .A1(n1390), .A2(n1391), .ZN(n1385) );
NAND2_X1 U19460 ( .A1(n1392), .A2(n1393), .ZN(n1390) );
OR2_X1 U19461 ( .A1(n1319), .A2(ex_block_i_alu_i_shift_amt_compl_0), .ZN(n1393) );
NOR2_X1 U19462 ( .A1(n1315), .A2(n1396), .ZN(n1392) );
NAND2_X1 U19463 ( .A1(n19966), .A2(n16067), .ZN(n1132) );
NAND2_X1 U19464 ( .A1(n19966), .A2(n16065), .ZN(n1034) );
NAND2_X1 U19465 ( .A1(n19966), .A2(n16064), .ZN(n996) );
NAND2_X1 U19466 ( .A1(n19966), .A2(n16063), .ZN(n957) );
NAND2_X1 U19467 ( .A1(n19966), .A2(n16062), .ZN(n918) );
NAND2_X1 U19468 ( .A1(n19966), .A2(n16061), .ZN(n837) );
NAND2_X1 U19469 ( .A1(n19966), .A2(n16060), .ZN(n798) );
NAND2_X1 U19470 ( .A1(n19966), .A2(n16059), .ZN(n760) );
NAND2_X1 U19471 ( .A1(n19966), .A2(n16058), .ZN(n723) );
NAND2_X1 U19472 ( .A1(n19966), .A2(n16072), .ZN(n39) );
NAND2_X1 U19473 ( .A1(n19966), .A2(n16071), .ZN(n1288) );
NAND2_X1 U19474 ( .A1(n19966), .A2(n16070), .ZN(n1249) );
NAND2_X1 U19475 ( .A1(n19966), .A2(n16069), .ZN(n1210) );
NAND2_X1 U19476 ( .A1(n19966), .A2(n16068), .ZN(n1171) );
NAND2_X1 U19477 ( .A1(n16346), .A2(n16066), .ZN(n1093) );
NAND2_X1 U19478 ( .A1(n1351), .A2(n1039), .ZN(n363) );
NOR2_X1 U19479 ( .A1(n1304), .A2(n33), .ZN(n1351) );
NAND2_X1 U19480 ( .A1(n16346), .A2(n16075), .ZN(n190) );
NAND2_X1 U19481 ( .A1(n16346), .A2(n16074), .ZN(n142) );
NAND2_X1 U19482 ( .A1(n16346), .A2(n16073), .ZN(n99) );
INV_X1 U19483 ( .A(n5128), .ZN(n20893) );
NAND2_X1 U19484 ( .A1(n1349), .A2(n1039), .ZN(n44) );
NOR2_X1 U19485 ( .A1(n1305), .A2(n33), .ZN(n1349) );
INV_X1 U19486 ( .A(n107), .ZN(n20718) );
INV_X1 U19487 ( .A(n51), .ZN(n20714) );
INV_X1 U19488 ( .A(n1295), .ZN(n20710) );
INV_X1 U19489 ( .A(n1217), .ZN(n20702) );
INV_X1 U19490 ( .A(n1178), .ZN(n20698) );
INV_X1 U19491 ( .A(n1139), .ZN(n20694) );
INV_X1 U19492 ( .A(n965), .ZN(n20645) );
INV_X1 U19493 ( .A(n926), .ZN(n20607) );
INV_X1 U19494 ( .A(n845), .ZN(n20567) );
INV_X1 U19495 ( .A(n768), .ZN(n20487) );
INV_X1 U19496 ( .A(n730), .ZN(n20447) );
INV_X1 U19497 ( .A(n693), .ZN(n20407) );
INV_X1 U19498 ( .A(n655), .ZN(n20368) );
INV_X1 U19499 ( .A(n615), .ZN(n20329) );
INV_X1 U19500 ( .A(n575), .ZN(n20290) );
INV_X1 U19501 ( .A(n535), .ZN(n20251) );
INV_X1 U19502 ( .A(n495), .ZN(n20213) );
INV_X1 U19503 ( .A(n806), .ZN(n20527) );
INV_X1 U19504 ( .A(n1003), .ZN(n20679) );
NAND2_X1 U19505 ( .A1(n7692), .A2(n7693), .ZN(n7691) );
NAND2_X1 U19506 ( .A1(n20993), .A2(n10304), .ZN(n10303) );
NAND2_X1 U19507 ( .A1(n20982), .A2(n5189), .ZN(n10304) );
INV_X1 U19508 ( .A(n5167), .ZN(n20982) );
NAND2_X1 U19509 ( .A1(n19967), .A2(n1354), .ZN(n1353) );
NAND2_X1 U19510 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
NOR2_X1 U19511 ( .A1(n1362), .A2(n1363), .ZN(n1355) );
NOR2_X1 U19512 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
OR2_X1 U19513 ( .A1(n20014), .A2(n1058), .ZN(n1057) );
AND2_X1 U19514 ( .A1(n16129), .A2(n7653), .ZN(n7698) );
NOR2_X1 U19515 ( .A1(n20961), .A2(n21002), .ZN(n6227) );
NAND2_X1 U19516 ( .A1(n7019), .A2(n7630), .ZN(n6793) );
NAND2_X1 U19517 ( .A1(n7030), .A2(n7019), .ZN(n6796) );
NOR2_X1 U19518 ( .A1(n15894), .A2(n7025), .ZN(n7030) );
NAND2_X1 U19519 ( .A1(n5088), .A2(n4959), .ZN(n5272) );
NAND2_X1 U19520 ( .A1(n15793), .A2(crash_dump_o_65_), .ZN(n2756) );
NOR2_X1 U19521 ( .A1(n1326), .A2(n1305), .ZN(n71) );
NAND2_X1 U19522 ( .A1(n4958), .A2(n5087), .ZN(n5586) );
NAND2_X1 U19523 ( .A1(n4958), .A2(n5088), .ZN(n5274) );
BUF_X1 U19524 ( .A(n2897), .Z(n16445) );
NAND2_X1 U19525 ( .A1(n5091), .A2(n20912), .ZN(n5090) );
AND2_X1 U19526 ( .A1(n10022), .A2(n15924), .ZN(n5908) );
BUF_X1 U19527 ( .A(n8557), .Z(n16376) );
BUF_X1 U19528 ( .A(n3129), .Z(n16436) );
BUF_X1 U19529 ( .A(n3262), .Z(n16434) );
NOR2_X1 U19530 ( .A1(n5550), .A2(n15887), .ZN(n4425) );
NAND2_X1 U19531 ( .A1(n5669), .A2(n20962), .ZN(n5374) );
NOR2_X1 U19532 ( .A1(n1435), .A2(n1431), .ZN(n5669) );
NOR2_X1 U19533 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N218), .A2(n11256), .ZN(n5011) );
NAND2_X1 U19534 ( .A1(crash_dump_o_65_), .A2(n15803), .ZN(n2164) );
NOR2_X1 U19535 ( .A1(n15815), .A2(n15918), .ZN(n10287) );
NOR2_X1 U19536 ( .A1(n6540), .A2(n15858), .ZN(n1564) );
NOR2_X1 U19537 ( .A1(n15925), .A2(n15825), .ZN(n1579) );
NOR2_X1 U19538 ( .A1(n1564), .A2(n1590), .ZN(n1565) );
NAND2_X1 U19539 ( .A1(n11255), .A2(n11254), .ZN(n22100) );
NAND2_X1 U19540 ( .A1(n4050), .A2(n4051), .ZN(n3777) );
NAND2_X1 U19541 ( .A1(n20985), .A2(n15813), .ZN(n4050) );
NOR2_X1 U19542 ( .A1(n15817), .A2(n15913), .ZN(n5245) );
NOR2_X1 U19543 ( .A1(n7041), .A2(n15919), .ZN(n7580) );
NAND2_X1 U19544 ( .A1(n9302), .A2(n9303), .ZN(n6896) );
NAND2_X1 U19545 ( .A1(n9304), .A2(n20527), .ZN(n9303) );
NAND2_X1 U19546 ( .A1(n806), .A2(n5268), .ZN(n9302) );
NOR2_X1 U19547 ( .A1(n19770), .A2(n16376), .ZN(n9304) );
NAND2_X1 U19548 ( .A1(n9514), .A2(n9515), .ZN(n6943) );
NAND2_X1 U19549 ( .A1(n9516), .A2(n20679), .ZN(n9515) );
NAND2_X1 U19550 ( .A1(n1003), .A2(n5268), .ZN(n9514) );
NOR2_X1 U19551 ( .A1(n19778), .A2(n16376), .ZN(n9516) );
NOR2_X1 U19552 ( .A1(n5112), .A2(n1444), .ZN(n1576) );
INV_X1 U19553 ( .A(n1040), .ZN(n21014) );
NAND2_X1 U19554 ( .A1(n3561), .A2(n3562), .ZN(n3126) );
NOR2_X1 U19555 ( .A1(n3563), .A2(n3564), .ZN(n3562) );
NOR2_X1 U19556 ( .A1(n3569), .A2(n3570), .ZN(n3561) );
NOR2_X1 U19557 ( .A1(n3565), .A2(n15812), .ZN(n3564) );
NAND2_X1 U19558 ( .A1(n19942), .A2(n2727), .ZN(n2058) );
NAND2_X1 U19559 ( .A1(n10353), .A2(n10354), .ZN(n1435) );
NOR2_X1 U19560 ( .A1(n10397), .A2(n10398), .ZN(n10353) );
NOR2_X1 U19561 ( .A1(n10355), .A2(n10356), .ZN(n10354) );
NAND2_X1 U19562 ( .A1(n10399), .A2(n10400), .ZN(n10397) );
NAND2_X1 U19563 ( .A1(n9712), .A2(n9713), .ZN(n7068) );
NAND2_X1 U19564 ( .A1(n9714), .A2(n20702), .ZN(n9713) );
NAND2_X1 U19565 ( .A1(n1217), .A2(n5268), .ZN(n9712) );
NOR2_X1 U19566 ( .A1(n19788), .A2(n8557), .ZN(n9714) );
NAND2_X1 U19567 ( .A1(n9752), .A2(n9753), .ZN(n7069) );
NAND2_X1 U19568 ( .A1(n9754), .A2(n20706), .ZN(n9753) );
NAND2_X1 U19569 ( .A1(n1258), .A2(n5268), .ZN(n9752) );
INV_X1 U19570 ( .A(n1258), .ZN(n20706) );
NAND2_X1 U19571 ( .A1(n9056), .A2(n9057), .ZN(n6842) );
NAND2_X1 U19572 ( .A1(n9058), .A2(n20290), .ZN(n9057) );
NAND2_X1 U19573 ( .A1(n575), .A2(n16418), .ZN(n9056) );
NOR2_X1 U19574 ( .A1(n19758), .A2(n16376), .ZN(n9058) );
NAND2_X1 U19575 ( .A1(n9097), .A2(n9098), .ZN(n6851) );
NAND2_X1 U19576 ( .A1(n9099), .A2(n20329), .ZN(n9098) );
NAND2_X1 U19577 ( .A1(n615), .A2(n16418), .ZN(n9097) );
NOR2_X1 U19578 ( .A1(n19760), .A2(n16376), .ZN(n9099) );
NAND2_X1 U19579 ( .A1(n9138), .A2(n9139), .ZN(n6860) );
NAND2_X1 U19580 ( .A1(n9140), .A2(n20368), .ZN(n9139) );
NAND2_X1 U19581 ( .A1(n655), .A2(n16418), .ZN(n9138) );
NOR2_X1 U19582 ( .A1(n19762), .A2(n16376), .ZN(n9140) );
NAND2_X1 U19583 ( .A1(n9179), .A2(n9180), .ZN(n6869) );
NAND2_X1 U19584 ( .A1(n9181), .A2(n20407), .ZN(n9180) );
NAND2_X1 U19585 ( .A1(n693), .A2(n5268), .ZN(n9179) );
NOR2_X1 U19586 ( .A1(n19764), .A2(n16376), .ZN(n9181) );
NAND2_X1 U19587 ( .A1(n9220), .A2(n9221), .ZN(n6878) );
NAND2_X1 U19588 ( .A1(n9222), .A2(n20447), .ZN(n9221) );
NAND2_X1 U19589 ( .A1(n730), .A2(n16418), .ZN(n9220) );
NOR2_X1 U19590 ( .A1(n19766), .A2(n16376), .ZN(n9222) );
NAND2_X1 U19591 ( .A1(n9261), .A2(n9262), .ZN(n6887) );
NAND2_X1 U19592 ( .A1(n9263), .A2(n20487), .ZN(n9262) );
NAND2_X1 U19593 ( .A1(n768), .A2(n5268), .ZN(n9261) );
NOR2_X1 U19594 ( .A1(n19768), .A2(n16376), .ZN(n9263) );
NAND2_X1 U19595 ( .A1(n9345), .A2(n9346), .ZN(n6905) );
NAND2_X1 U19596 ( .A1(n9347), .A2(n20567), .ZN(n9346) );
NAND2_X1 U19597 ( .A1(n845), .A2(n16418), .ZN(n9345) );
NOR2_X1 U19598 ( .A1(n19772), .A2(n16376), .ZN(n9347) );
NAND2_X1 U19599 ( .A1(n9432), .A2(n9433), .ZN(n6925) );
NAND2_X1 U19600 ( .A1(n9434), .A2(n20607), .ZN(n9433) );
NAND2_X1 U19601 ( .A1(n926), .A2(n5268), .ZN(n9432) );
NOR2_X1 U19602 ( .A1(n19774), .A2(n16376), .ZN(n9434) );
NAND2_X1 U19603 ( .A1(n9473), .A2(n9474), .ZN(n6934) );
NAND2_X1 U19604 ( .A1(n9475), .A2(n20645), .ZN(n9474) );
NAND2_X1 U19605 ( .A1(n965), .A2(n16418), .ZN(n9473) );
NOR2_X1 U19606 ( .A1(n19776), .A2(n8557), .ZN(n9475) );
NAND2_X1 U19607 ( .A1(n9558), .A2(n9559), .ZN(n6952) );
NAND2_X1 U19608 ( .A1(n9560), .A2(n20686), .ZN(n9559) );
NAND2_X1 U19609 ( .A1(n1046), .A2(n5268), .ZN(n9558) );
INV_X1 U19610 ( .A(n1046), .ZN(n20686) );
NAND2_X1 U19611 ( .A1(n9848), .A2(n9849), .ZN(n7203) );
NAND2_X1 U19612 ( .A1(n9850), .A2(n20751), .ZN(n9849) );
NAND2_X1 U19613 ( .A1(n466), .A2(n5268), .ZN(n9848) );
NOR2_X1 U19614 ( .A1(n19808), .A2(n16376), .ZN(n9850) );
NAND2_X1 U19615 ( .A1(n9015), .A2(n9016), .ZN(n6833) );
NAND2_X1 U19616 ( .A1(n9017), .A2(n20251), .ZN(n9016) );
NAND2_X1 U19617 ( .A1(n535), .A2(n16418), .ZN(n9015) );
NOR2_X1 U19618 ( .A1(n19756), .A2(n16376), .ZN(n9017) );
NAND2_X1 U19619 ( .A1(n8974), .A2(n8975), .ZN(n6824) );
NAND2_X1 U19620 ( .A1(n8976), .A2(n20213), .ZN(n8975) );
NAND2_X1 U19621 ( .A1(n495), .A2(n16418), .ZN(n8974) );
NOR2_X1 U19622 ( .A1(n19754), .A2(n16376), .ZN(n8976) );
NAND2_X1 U19623 ( .A1(n8927), .A2(n8928), .ZN(n6803) );
NAND2_X1 U19624 ( .A1(n8929), .A2(n20175), .ZN(n8928) );
NAND2_X1 U19625 ( .A1(n414), .A2(n16418), .ZN(n8927) );
INV_X1 U19626 ( .A(n414), .ZN(n20175) );
NAND2_X1 U19627 ( .A1(n10526), .A2(n10527), .ZN(n10051) );
NOR2_X1 U19628 ( .A1(n20979), .A2(n10529), .ZN(n10527) );
NOR2_X1 U19629 ( .A1(n10156), .A2(n9968), .ZN(n10526) );
INV_X1 U19630 ( .A(n10150), .ZN(n20979) );
NOR2_X1 U19631 ( .A1(crash_dump_o_65_), .A2(n3050), .ZN(n1447) );
INV_X1 U19632 ( .A(n7722), .ZN(n20988) );
NOR2_X1 U19633 ( .A1(n2042), .A2(n2456), .ZN(n2539) );
NOR2_X1 U19634 ( .A1(n15879), .A2(n15805), .ZN(n10367) );
NOR2_X1 U19635 ( .A1(n15860), .A2(n10193), .ZN(n10204) );
NAND2_X1 U19636 ( .A1(n19905), .A2(n2042), .ZN(n2409) );
INV_X1 U19637 ( .A(n1444), .ZN(n20990) );
NOR2_X1 U19638 ( .A1(n15915), .A2(n15819), .ZN(n10461) );
INV_X1 U19639 ( .A(n1575), .ZN(n20993) );
NAND2_X1 U19640 ( .A1(n10535), .A2(n20994), .ZN(n10156) );
AND2_X1 U19641 ( .A1(n10144), .A2(n10143), .ZN(n10535) );
NAND2_X1 U19642 ( .A1(n21004), .A2(n15877), .ZN(n4431) );
NAND2_X1 U19643 ( .A1(n20922), .A2(n5671), .ZN(n4940) );
NAND2_X1 U19644 ( .A1(n9600), .A2(n9601), .ZN(n7237) );
NAND2_X1 U19645 ( .A1(n9602), .A2(n20690), .ZN(n9601) );
NAND2_X1 U19646 ( .A1(n1102), .A2(n5268), .ZN(n9600) );
INV_X1 U19647 ( .A(n1102), .ZN(n20690) );
NAND2_X1 U19648 ( .A1(n9675), .A2(n9676), .ZN(n7243) );
NAND2_X1 U19649 ( .A1(n9677), .A2(n20698), .ZN(n9676) );
NAND2_X1 U19650 ( .A1(n1178), .A2(n5268), .ZN(n9675) );
NOR2_X1 U19651 ( .A1(n19786), .A2(n16376), .ZN(n9677) );
NAND2_X1 U19652 ( .A1(n8649), .A2(n8650), .ZN(n7185) );
NAND2_X1 U19653 ( .A1(n8651), .A2(n20723), .ZN(n8650) );
NAND2_X1 U19654 ( .A1(n170), .A2(n16418), .ZN(n8649) );
NOR2_X1 U19655 ( .A1(n19798), .A2(n8557), .ZN(n8651) );
NAND2_X1 U19656 ( .A1(n8892), .A2(n8893), .ZN(n6792) );
NAND2_X1 U19657 ( .A1(n8894), .A2(n20136), .ZN(n8893) );
NAND2_X1 U19658 ( .A1(n5268), .A2(n5799), .ZN(n8892) );
NOR2_X1 U19659 ( .A1(n19750), .A2(n8557), .ZN(n8894) );
INV_X1 U19660 ( .A(n2042), .ZN(n19914) );
NOR2_X1 U19661 ( .A1(n1580), .A2(n1581), .ZN(n1525) );
NOR2_X1 U19662 ( .A1(n1553), .A2(n1528), .ZN(n1531) );
NAND2_X1 U19663 ( .A1(n20986), .A2(n5182), .ZN(n5147) );
NAND2_X1 U19664 ( .A1(n1689), .A2(n1690), .ZN(n1606) );
NOR2_X1 U19665 ( .A1(n1693), .A2(n1694), .ZN(n1689) );
NOR2_X1 U19666 ( .A1(n1538), .A2(n1691), .ZN(n1690) );
NOR2_X1 U19667 ( .A1(n1695), .A2(n19965), .ZN(n1694) );
NAND2_X1 U19668 ( .A1(n9965), .A2(n20948), .ZN(n8819) );
NOR2_X1 U19669 ( .A1(n20949), .A2(n9968), .ZN(n9965) );
NAND2_X1 U19670 ( .A1(n2851), .A2(n19910), .ZN(n2715) );
NOR2_X1 U19671 ( .A1(n19907), .A2(n2440), .ZN(n2851) );
NAND2_X1 U19672 ( .A1(n4939), .A2(n10292), .ZN(n5091) );
NAND2_X1 U19673 ( .A1(n10293), .A2(n20971), .ZN(n10292) );
INV_X1 U19674 ( .A(n5583), .ZN(n20971) );
NOR2_X1 U19675 ( .A1(n10185), .A2(n5580), .ZN(n10293) );
NAND2_X1 U19676 ( .A1(n2437), .A2(n2035), .ZN(n2410) );
NAND2_X1 U19677 ( .A1(n10205), .A2(n10206), .ZN(n1395) );
NOR2_X1 U19678 ( .A1(n10214), .A2(n10197), .ZN(n10205) );
NOR2_X1 U19679 ( .A1(n10207), .A2(n10208), .ZN(n10206) );
NOR2_X1 U19680 ( .A1(n10203), .A2(n10188), .ZN(n10214) );
AND2_X1 U19681 ( .A1(n20906), .A2(n5665), .ZN(n5651) );
NAND2_X1 U19682 ( .A1(n5556), .A2(n4927), .ZN(n5665) );
NAND2_X1 U19683 ( .A1(n10176), .A2(n10177), .ZN(n6231) );
NOR2_X1 U19684 ( .A1(n10196), .A2(n10197), .ZN(n10176) );
NOR2_X1 U19685 ( .A1(n10178), .A2(n10179), .ZN(n10177) );
NOR2_X1 U19686 ( .A1(n10198), .A2(n10182), .ZN(n10196) );
NOR2_X1 U19687 ( .A1(n2042), .A2(n19927), .ZN(n2702) );
INV_X1 U19688 ( .A(n1507), .ZN(n19963) );
NAND2_X1 U19689 ( .A1(n9638), .A2(n9639), .ZN(n7240) );
NAND2_X1 U19690 ( .A1(n9640), .A2(n20694), .ZN(n9639) );
NAND2_X1 U19691 ( .A1(n1139), .A2(n5268), .ZN(n9638) );
NOR2_X1 U19692 ( .A1(n19784), .A2(n8557), .ZN(n9640) );
NAND2_X1 U19693 ( .A1(n9800), .A2(n9801), .ZN(n7250) );
NAND2_X1 U19694 ( .A1(n9802), .A2(n20710), .ZN(n9801) );
NAND2_X1 U19695 ( .A1(n1295), .A2(n5268), .ZN(n9800) );
NOR2_X1 U19696 ( .A1(n19792), .A2(n16376), .ZN(n9802) );
NAND2_X1 U19697 ( .A1(n8553), .A2(n8554), .ZN(n7179) );
NAND2_X1 U19698 ( .A1(n8555), .A2(n20714), .ZN(n8554) );
NAND2_X1 U19699 ( .A1(n51), .A2(n16418), .ZN(n8553) );
NOR2_X1 U19700 ( .A1(n19794), .A2(n8557), .ZN(n8555) );
NAND2_X1 U19701 ( .A1(n8606), .A2(n8607), .ZN(n7182) );
NAND2_X1 U19702 ( .A1(n8608), .A2(n20718), .ZN(n8607) );
NAND2_X1 U19703 ( .A1(n107), .A2(n16418), .ZN(n8606) );
NOR2_X1 U19704 ( .A1(n19796), .A2(n8557), .ZN(n8608) );
NAND2_X1 U19705 ( .A1(n8697), .A2(n8698), .ZN(n7188) );
NAND2_X1 U19706 ( .A1(n8699), .A2(n20729), .ZN(n8698) );
NAND2_X1 U19707 ( .A1(n213), .A2(n16418), .ZN(n8697) );
NOR2_X1 U19708 ( .A1(n19800), .A2(n8557), .ZN(n8699) );
NAND2_X1 U19709 ( .A1(n9894), .A2(n9895), .ZN(n7253) );
NAND2_X1 U19710 ( .A1(n9896), .A2(n20759), .ZN(n9895) );
NAND2_X1 U19711 ( .A1(n1391), .A2(n16418), .ZN(n9894) );
NOR2_X1 U19712 ( .A1(n19812), .A2(n16376), .ZN(n9896) );
NAND2_X1 U19713 ( .A1(n8734), .A2(n8735), .ZN(n7191) );
NAND2_X1 U19714 ( .A1(n8736), .A2(n20734), .ZN(n8735) );
NAND2_X1 U19715 ( .A1(n240), .A2(n16418), .ZN(n8734) );
INV_X1 U19716 ( .A(n240), .ZN(n20734) );
INV_X1 U19717 ( .A(n3042), .ZN(n19885) );
NOR2_X1 U19718 ( .A1(n1549), .A2(n1571), .ZN(n1553) );
NOR2_X1 U19719 ( .A1(n21005), .A2(n4431), .ZN(n5547) );
INV_X1 U19720 ( .A(n5542), .ZN(n21005) );
NOR2_X1 U19721 ( .A1(n1564), .A2(n20934), .ZN(n6526) );
INV_X1 U19722 ( .A(n6525), .ZN(n20934) );
NAND2_X1 U19723 ( .A1(n15923), .A2(n15822), .ZN(n1058) );
NOR2_X1 U19724 ( .A1(n5198), .A2(n5221), .ZN(n5184) );
NOR2_X1 U19725 ( .A1(n1575), .A2(n1576), .ZN(n1520) );
NOR2_X1 U19726 ( .A1(n5127), .A2(n5209), .ZN(n5183) );
NAND2_X1 U19727 ( .A1(n5210), .A2(n5151), .ZN(n5209) );
NOR2_X1 U19728 ( .A1(n10274), .A2(n1435), .ZN(data_we_o) );
INV_X1 U19729 ( .A(n4939), .ZN(n20962) );
NOR2_X1 U19730 ( .A1(n22094), .A2(n22089), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_18) );
NOR2_X1 U19731 ( .A1(n22094), .A2(n22090), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_19) );
NOR2_X1 U19732 ( .A1(n22095), .A2(n22089), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_20) );
NOR2_X1 U19733 ( .A1(n22095), .A2(n22090), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_21) );
NOR2_X1 U19734 ( .A1(n22094), .A2(n22092), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_26) );
NOR2_X1 U19735 ( .A1(n22094), .A2(n22093), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_27) );
NOR2_X1 U19736 ( .A1(n22095), .A2(n22092), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_28) );
NOR2_X1 U19737 ( .A1(n22095), .A2(n22093), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_29) );
NOR2_X1 U19738 ( .A1(n22097), .A2(n22093), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_31) );
NOR2_X1 U19739 ( .A1(n22097), .A2(n22089), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_22) );
NOR2_X1 U19740 ( .A1(n22097), .A2(n22090), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_23) );
NOR2_X1 U19741 ( .A1(n22097), .A2(n22092), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_30) );
NAND2_X1 U19742 ( .A1(n16451), .A2(n2042), .ZN(n2441) );
NOR2_X1 U19743 ( .A1(n22100), .A2(n22090), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_17) );
NOR2_X1 U19744 ( .A1(n22100), .A2(n22093), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_25) );
NOR2_X1 U19745 ( .A1(n10172), .A2(n10182), .ZN(n10166) );
NOR2_X1 U19746 ( .A1(n10449), .A2(n5138), .ZN(n6701) );
OR2_X1 U19747 ( .A1(n5182), .A2(n4056), .ZN(n10449) );
NOR2_X1 U19748 ( .A1(n5167), .A2(n5189), .ZN(n5153) );
INV_X1 U19749 ( .A(n2136), .ZN(n19929) );
INV_X1 U19750 ( .A(n2440), .ZN(n19912) );
NOR2_X1 U19751 ( .A1(n10224), .A2(n10204), .ZN(n10103) );
NOR2_X1 U19752 ( .A1(n20970), .A2(n15860), .ZN(n10224) );
INV_X1 U19753 ( .A(n5010), .ZN(n21007) );
NOR2_X1 U19754 ( .A1(n15810), .A2(n15859), .ZN(n10169) );
NOR2_X1 U19755 ( .A1(n5269), .A2(n10438), .ZN(n10425) );
NOR2_X1 U19756 ( .A1(n15793), .A2(n2753), .ZN(n2746) );
NAND2_X1 U19757 ( .A1(n3699), .A2(n3700), .ZN(n1446) );
NOR2_X1 U19758 ( .A1(n20895), .A2(n3702), .ZN(n3700) );
NOR2_X1 U19759 ( .A1(n15878), .A2(n15929), .ZN(n3699) );
NAND2_X1 U19760 ( .A1(n3703), .A2(n3704), .ZN(n3702) );
NAND2_X1 U19761 ( .A1(n10232), .A2(n20990), .ZN(n6306) );
NOR2_X1 U19762 ( .A1(n10233), .A2(n10234), .ZN(n10232) );
NAND2_X1 U19763 ( .A1(n16453), .A2(n2203), .ZN(n2024) );
AND2_X1 U19764 ( .A1(n5232), .A2(n5233), .ZN(n5198) );
NOR2_X1 U19765 ( .A1(n19986), .A2(n5253), .ZN(n5232) );
NOR2_X1 U19766 ( .A1(n15563), .A2(n20932), .ZN(n5233) );
INV_X1 U19767 ( .A(n5116), .ZN(n19986) );
NOR2_X1 U19768 ( .A1(n15924), .A2(n15824), .ZN(n10390) );
INV_X1 U19769 ( .A(n2043), .ZN(n19934) );
NOR2_X1 U19770 ( .A1(n2136), .A2(n2018), .ZN(n2773) );
INV_X1 U19771 ( .A(n4056), .ZN(n20986) );
NOR2_X1 U19772 ( .A1(n5556), .A2(n15877), .ZN(n5540) );
INV_X1 U19773 ( .A(n4435), .ZN(n20110) );
NOR2_X1 U19774 ( .A1(n2782), .A2(n19908), .ZN(n2893) );
NOR2_X1 U19775 ( .A1(n2782), .A2(n19911), .ZN(n2877) );
NOR2_X1 U19776 ( .A1(n2782), .A2(n19920), .ZN(n2843) );
NOR2_X1 U19777 ( .A1(n2782), .A2(n19913), .ZN(n2885) );
NOR2_X1 U19778 ( .A1(n2782), .A2(n19928), .ZN(n2804) );
NOR2_X1 U19779 ( .A1(n2782), .A2(n19915), .ZN(n2849) );
NOR2_X1 U19780 ( .A1(n2782), .A2(n19924), .ZN(n2836) );
NOR2_X1 U19781 ( .A1(n2782), .A2(n19926), .ZN(n2822) );
NOR2_X1 U19782 ( .A1(n2782), .A2(n19932), .ZN(n2781) );
NOR2_X1 U19783 ( .A1(n2782), .A2(n19935), .ZN(n2788) );
NOR2_X1 U19784 ( .A1(n2782), .A2(n19930), .ZN(n2812) );
NOR2_X1 U19785 ( .A1(n2782), .A2(n19933), .ZN(n2795) );
NOR2_X1 U19786 ( .A1(n2782), .A2(n19922), .ZN(n2828) );
NOR2_X1 U19787 ( .A1(n2782), .A2(n19918), .ZN(n2857) );
NAND2_X1 U19788 ( .A1(n19910), .A2(n2440), .ZN(n2522) );
INV_X1 U19789 ( .A(n2437), .ZN(n19910) );
NOR2_X1 U19790 ( .A1(n2042), .A2(n2470), .ZN(n2172) );
NOR2_X1 U19791 ( .A1(n15880), .A2(n5911), .ZN(n6178) );
NOR2_X1 U19792 ( .A1(n15881), .A2(n5911), .ZN(n6164) );
NOR2_X1 U19793 ( .A1(n15882), .A2(n5911), .ZN(n6150) );
NOR2_X1 U19794 ( .A1(n15883), .A2(n5911), .ZN(n6137) );
NOR2_X1 U19795 ( .A1(n15861), .A2(n5911), .ZN(n6124) );
NOR2_X1 U19796 ( .A1(n15862), .A2(n5911), .ZN(n6110) );
NOR2_X1 U19797 ( .A1(n15863), .A2(n5911), .ZN(n6096) );
NOR2_X1 U19798 ( .A1(n15864), .A2(n5911), .ZN(n6070) );
NOR2_X1 U19799 ( .A1(n15865), .A2(n5911), .ZN(n6056) );
NOR2_X1 U19800 ( .A1(n15866), .A2(n5911), .ZN(n6042) );
NOR2_X1 U19801 ( .A1(n15867), .A2(n5911), .ZN(n6028) );
NOR2_X1 U19802 ( .A1(n15868), .A2(n5911), .ZN(n6014) );
NOR2_X1 U19803 ( .A1(n15869), .A2(n5911), .ZN(n6000) );
NOR2_X1 U19804 ( .A1(n15870), .A2(n5911), .ZN(n5986) );
NOR2_X1 U19805 ( .A1(n15871), .A2(n5911), .ZN(n5972) );
NOR2_X1 U19806 ( .A1(n15872), .A2(n5911), .ZN(n5958) );
NOR2_X1 U19807 ( .A1(n15873), .A2(n5911), .ZN(n5944) );
NOR2_X1 U19808 ( .A1(n15874), .A2(n5911), .ZN(n5920) );
NOR2_X1 U19809 ( .A1(n15875), .A2(n5911), .ZN(n5900) );
NAND2_X1 U19810 ( .A1(n19909), .A2(n2042), .ZN(n2303) );
NAND2_X1 U19811 ( .A1(n22086), .A2(n11256), .ZN(n22099) );
NAND2_X1 U19812 ( .A1(n5687), .A2(n5709), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_18) );
NAND2_X1 U19813 ( .A1(n16412), .A2(n15863), .ZN(n5709) );
NAND2_X1 U19814 ( .A1(n5687), .A2(n5708), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_19) );
NAND2_X1 U19815 ( .A1(n16412), .A2(n15864), .ZN(n5708) );
NAND2_X1 U19816 ( .A1(n5687), .A2(n5705), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_20) );
NAND2_X1 U19817 ( .A1(n16412), .A2(n15865), .ZN(n5705) );
NAND2_X1 U19818 ( .A1(n5687), .A2(n5704), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_21) );
NAND2_X1 U19819 ( .A1(n16412), .A2(n15866), .ZN(n5704) );
NAND2_X1 U19820 ( .A1(n5687), .A2(n5703), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_22) );
NAND2_X1 U19821 ( .A1(n16412), .A2(n15867), .ZN(n5703) );
NAND2_X1 U19822 ( .A1(n5687), .A2(n5702), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_23) );
NAND2_X1 U19823 ( .A1(n16412), .A2(n15868), .ZN(n5702) );
NAND2_X1 U19824 ( .A1(n5687), .A2(n5701), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_24) );
NAND2_X1 U19825 ( .A1(n16412), .A2(n15869), .ZN(n5701) );
NAND2_X1 U19826 ( .A1(n5687), .A2(n5700), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_25) );
NAND2_X1 U19827 ( .A1(n16412), .A2(n15870), .ZN(n5700) );
NAND2_X1 U19828 ( .A1(n5687), .A2(n5699), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_26) );
NAND2_X1 U19829 ( .A1(n16412), .A2(n15871), .ZN(n5699) );
NAND2_X1 U19830 ( .A1(n5687), .A2(n5698), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_27) );
NAND2_X1 U19831 ( .A1(n16412), .A2(n15872), .ZN(n5698) );
NAND2_X1 U19832 ( .A1(n5687), .A2(n5697), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_28) );
NAND2_X1 U19833 ( .A1(n16412), .A2(n15873), .ZN(n5697) );
NAND2_X1 U19834 ( .A1(n5687), .A2(n5696), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_29) );
NAND2_X1 U19835 ( .A1(n16412), .A2(n15874), .ZN(n5696) );
NAND2_X1 U19836 ( .A1(n5687), .A2(n5693), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_30) );
NAND2_X1 U19837 ( .A1(n16411), .A2(n15875), .ZN(n5693) );
NAND2_X1 U19838 ( .A1(n5687), .A2(n5692), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_31) );
NAND2_X1 U19839 ( .A1(n16411), .A2(n15891), .ZN(n5692) );
NAND2_X1 U19840 ( .A1(n5687), .A2(n5690), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_32) );
NAND2_X1 U19841 ( .A1(n16411), .A2(n15930), .ZN(n5690) );
NAND2_X1 U19842 ( .A1(n22088), .A2(n11256), .ZN(n22096) );
INV_X1 U19843 ( .A(n1581), .ZN(n20996) );
NAND2_X1 U19844 ( .A1(n22087), .A2(n11256), .ZN(n22089) );
NAND2_X1 U19845 ( .A1(n22091), .A2(n11256), .ZN(n22092) );
NAND2_X1 U19846 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N218), .A2(n11256), .ZN(n4998) );
INV_X1 U19847 ( .A(n4996), .ZN(n21006) );
NAND2_X1 U19848 ( .A1(n10218), .A2(n10219), .ZN(n6234) );
NOR2_X1 U19849 ( .A1(n10235), .A2(n10148), .ZN(n10218) );
NOR2_X1 U19850 ( .A1(n10220), .A2(n10221), .ZN(n10219) );
NOR2_X1 U19851 ( .A1(n10249), .A2(n10185), .ZN(n10235) );
NAND2_X1 U19852 ( .A1(n2204), .A2(n2665), .ZN(n2566) );
NAND2_X1 U19853 ( .A1(n2141), .A2(n2042), .ZN(n2665) );
NAND2_X1 U19854 ( .A1(n15921), .A2(n15820), .ZN(n1597) );
NAND2_X1 U19855 ( .A1(n2773), .A2(n2774), .ZN(n2456) );
NOR2_X1 U19856 ( .A1(n2203), .A2(n2775), .ZN(n2774) );
NAND2_X1 U19857 ( .A1(n19934), .A2(n19931), .ZN(n2775) );
NAND2_X1 U19858 ( .A1(n10075), .A2(n10076), .ZN(n5222) );
NOR2_X1 U19859 ( .A1(n5108), .A2(n10268), .ZN(n10075) );
NOR2_X1 U19860 ( .A1(n15773), .A2(n10077), .ZN(n10076) );
NOR2_X1 U19861 ( .A1(n1431), .A2(n5115), .ZN(n10268) );
NAND2_X1 U19862 ( .A1(n1518), .A2(n10536), .ZN(n1687) );
NAND2_X1 U19863 ( .A1(n20995), .A2(n15916), .ZN(n10536) );
NAND2_X1 U19864 ( .A1(n9971), .A2(n9972), .ZN(n7084) );
AND2_X1 U19865 ( .A1(n9973), .A2(n8430), .ZN(n9972) );
NOR2_X1 U19866 ( .A1(n1431), .A2(n5222), .ZN(n9971) );
NAND2_X1 U19867 ( .A1(n10410), .A2(n10411), .ZN(n1596) );
NOR2_X1 U19868 ( .A1(n15876), .A2(n15804), .ZN(n10410) );
NOR2_X1 U19869 ( .A1(n15895), .A2(n10377), .ZN(n10411) );
NOR2_X1 U19870 ( .A1(n22097), .A2(n22096), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_6) );
NAND2_X1 U19871 ( .A1(n15908), .A2(n15799), .ZN(n10150) );
NAND2_X1 U19872 ( .A1(n5251), .A2(n20932), .ZN(n5173) );
NOR2_X1 U19873 ( .A1(n22100), .A2(n22098), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_1) );
NAND2_X1 U19874 ( .A1(n16450), .A2(n2591), .ZN(n2028) );
INV_X1 U19875 ( .A(n2426), .ZN(n19931) );
NAND2_X1 U19876 ( .A1(n2870), .A2(n19910), .ZN(n2349) );
NOR2_X1 U19877 ( .A1(n2035), .A2(n2440), .ZN(n2870) );
NOR2_X1 U19878 ( .A1(n15885), .A2(n6796), .ZN(n6926) );
NOR2_X1 U19879 ( .A1(n15806), .A2(n6796), .ZN(n6935) );
NOR2_X1 U19880 ( .A1(n15809), .A2(n6796), .ZN(n6953) );
NOR2_X1 U19881 ( .A1(n15889), .A2(n6796), .ZN(n6944) );
INV_X1 U19882 ( .A(n2169), .ZN(n16449) );
INV_X1 U19883 ( .A(n10185), .ZN(n20963) );
NOR2_X1 U19884 ( .A1(n22099), .A2(n22094), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_10) );
NOR2_X1 U19885 ( .A1(n22101), .A2(n22094), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_11) );
NOR2_X1 U19886 ( .A1(n22099), .A2(n22095), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_12) );
NOR2_X1 U19887 ( .A1(n22101), .A2(n22095), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_13) );
NOR2_X1 U19888 ( .A1(n22096), .A2(n22094), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_2) );
NOR2_X1 U19889 ( .A1(n22098), .A2(n22094), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_3) );
NOR2_X1 U19890 ( .A1(n22096), .A2(n22095), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_4) );
NOR2_X1 U19891 ( .A1(n22098), .A2(n22095), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_5) );
NOR2_X1 U19892 ( .A1(n22099), .A2(n22097), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_14) );
NOR2_X1 U19893 ( .A1(n22101), .A2(n22097), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_15) );
NOR2_X1 U19894 ( .A1(n22098), .A2(n22097), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_7) );
NOR2_X1 U19895 ( .A1(n22101), .A2(n22100), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_9) );
NOR2_X1 U19896 ( .A1(n5735), .A2(n4958), .ZN(n5736) );
NAND2_X1 U19897 ( .A1(n19899), .A2(n2042), .ZN(n2204) );
INV_X1 U19898 ( .A(n2170), .ZN(n16447) );
NOR2_X1 U19899 ( .A1(n10244), .A2(n10234), .ZN(n10516) );
NOR2_X1 U19900 ( .A1(n19945), .A2(n2782), .ZN(n2869) );
NAND2_X1 U19901 ( .A1(n20946), .A2(n15859), .ZN(n10203) );
NOR2_X1 U19902 ( .A1(n2170), .A2(n19935), .ZN(n2286) );
NAND2_X1 U19903 ( .A1(n10464), .A2(n15800), .ZN(n5120) );
NAND2_X1 U19904 ( .A1(n7722), .A2(n8127), .ZN(n8074) );
NAND2_X1 U19905 ( .A1(n19983), .A2(n16201), .ZN(n8127) );
NAND2_X1 U19906 ( .A1(n21000), .A2(n15877), .ZN(n4258) );
INV_X1 U19907 ( .A(n2782), .ZN(n20905) );
NOR2_X1 U19908 ( .A1(n16446), .A2(n19926), .ZN(n2167) );
NOR2_X1 U19909 ( .A1(n2170), .A2(n19920), .ZN(n2635) );
NOR2_X1 U19910 ( .A1(n16446), .A2(n19915), .ZN(n2578) );
NOR2_X1 U19911 ( .A1(n2170), .A2(n19918), .ZN(n2607) );
NOR2_X1 U19912 ( .A1(n16446), .A2(n19932), .ZN(n2229) );
NOR2_X1 U19913 ( .A1(n16446), .A2(n19946), .ZN(n2890) );
NOR2_X1 U19914 ( .A1(n16446), .A2(n19947), .ZN(n2874) );
NOR2_X1 U19915 ( .A1(n2170), .A2(n19951), .ZN(n2841) );
NOR2_X1 U19916 ( .A1(n16446), .A2(n19948), .ZN(n2882) );
NOR2_X1 U19917 ( .A1(n2170), .A2(n19955), .ZN(n2801) );
NOR2_X1 U19918 ( .A1(n16446), .A2(n19949), .ZN(n2847) );
NOR2_X1 U19919 ( .A1(n16446), .A2(n19953), .ZN(n2833) );
NOR2_X1 U19920 ( .A1(n16446), .A2(n19954), .ZN(n2820) );
NOR2_X1 U19921 ( .A1(n16446), .A2(n19957), .ZN(n2779) );
NOR2_X1 U19922 ( .A1(n2170), .A2(n19959), .ZN(n2786) );
NOR2_X1 U19923 ( .A1(n2170), .A2(n19956), .ZN(n2809) );
NOR2_X1 U19924 ( .A1(n16446), .A2(n19958), .ZN(n2792) );
NOR2_X1 U19925 ( .A1(n2170), .A2(n19952), .ZN(n2826) );
NOR2_X1 U19926 ( .A1(n2170), .A2(n19950), .ZN(n2855) );
NOR2_X1 U19927 ( .A1(n10433), .A2(rf_raddr_b_o_1_), .ZN(n5263) );
NOR2_X1 U19928 ( .A1(n2565), .A2(n19881), .ZN(n2562) );
NOR2_X1 U19929 ( .A1(n2566), .A2(n2567), .ZN(n2565) );
NAND2_X1 U19930 ( .A1(n2568), .A2(n2569), .ZN(n2567) );
NAND2_X1 U19931 ( .A1(n19904), .A2(n2570), .ZN(n2569) );
NOR2_X1 U19932 ( .A1(n2650), .A2(n19881), .ZN(n2645) );
NOR2_X1 U19933 ( .A1(n2566), .A2(n2651), .ZN(n2650) );
NAND2_X1 U19934 ( .A1(n2652), .A2(n2653), .ZN(n2651) );
NAND2_X1 U19935 ( .A1(n19904), .A2(n2644), .ZN(n2652) );
INV_X1 U19936 ( .A(n3019), .ZN(n19886) );
NAND2_X1 U19937 ( .A1(n5687), .A2(n5688), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_33) );
NAND2_X1 U19938 ( .A1(n16411), .A2(n15931), .ZN(n5688) );
NAND2_X1 U19939 ( .A1(n15922), .A2(n15823), .ZN(n5088) );
NOR2_X1 U19940 ( .A1(n2208), .A2(n2117), .ZN(n2206) );
NOR2_X1 U19941 ( .A1(n2209), .A2(n2210), .ZN(n2208) );
NAND2_X1 U19942 ( .A1(n2211), .A2(n2212), .ZN(n2210) );
NAND2_X1 U19943 ( .A1(n2214), .A2(n2215), .ZN(n2209) );
NOR2_X1 U19944 ( .A1(n2116), .A2(n2117), .ZN(n2114) );
NOR2_X1 U19945 ( .A1(n2118), .A2(n2119), .ZN(n2116) );
NAND2_X1 U19946 ( .A1(n2120), .A2(n2121), .ZN(n2119) );
NAND2_X1 U19947 ( .A1(n2125), .A2(n2126), .ZN(n2118) );
NOR2_X1 U19948 ( .A1(n19961), .A2(n2170), .ZN(n2867) );
NOR2_X1 U19949 ( .A1(n19960), .A2(n2170), .ZN(n2862) );
NOR2_X1 U19950 ( .A1(n2293), .A2(n2117), .ZN(n2292) );
NOR2_X1 U19951 ( .A1(n2294), .A2(n2295), .ZN(n2293) );
NOR2_X1 U19952 ( .A1(n2296), .A2(n2297), .ZN(n2295) );
NOR2_X1 U19953 ( .A1(n19943), .A2(crash_dump_o_65_), .ZN(n2294) );
NOR2_X1 U19954 ( .A1(n20853), .A2(n1297), .ZN(n8116) );
INV_X1 U19955 ( .A(n5550), .ZN(n21002) );
NOR2_X1 U19956 ( .A1(n3050), .A2(n2169), .ZN(n3584) );
NOR2_X1 U19957 ( .A1(n3050), .A2(n2170), .ZN(n3569) );
NOR2_X1 U19958 ( .A1(n19945), .A2(n16446), .ZN(n2329) );
NOR2_X1 U19959 ( .A1(n2035), .A2(n2036), .ZN(n2034) );
INV_X1 U19960 ( .A(n2103), .ZN(n19917) );
NAND2_X1 U19961 ( .A1(n20952), .A2(n15859), .ZN(n10172) );
INV_X1 U19962 ( .A(n2018), .ZN(n19927) );
NOR2_X1 U19963 ( .A1(n19949), .A2(n2166), .ZN(n2575) );
NOR2_X1 U19964 ( .A1(n19950), .A2(n2166), .ZN(n2604) );
NOR2_X1 U19965 ( .A1(n19954), .A2(n2166), .ZN(n2162) );
NOR2_X1 U19966 ( .A1(n19959), .A2(n2166), .ZN(n2283) );
NOR2_X1 U19967 ( .A1(n19961), .A2(n2166), .ZN(n2326) );
NOR2_X1 U19968 ( .A1(n16420), .A2(n15899), .ZN(n4403) );
NOR2_X1 U19969 ( .A1(n16420), .A2(n15900), .ZN(n4384) );
NOR2_X1 U19970 ( .A1(n16420), .A2(n15901), .ZN(n4365) );
NOR2_X1 U19971 ( .A1(n16420), .A2(n15902), .ZN(n4346) );
NOR2_X1 U19972 ( .A1(n16420), .A2(n15903), .ZN(n4327) );
NOR2_X1 U19973 ( .A1(n16420), .A2(n15904), .ZN(n4308) );
NOR2_X1 U19974 ( .A1(n16420), .A2(n15905), .ZN(n4285) );
NAND2_X1 U19975 ( .A1(n20933), .A2(n15907), .ZN(n5249) );
NAND2_X1 U19976 ( .A1(n20994), .A2(n10513), .ZN(n10493) );
NAND2_X1 U19977 ( .A1(n10514), .A2(n10145), .ZN(n10513) );
NOR2_X1 U19978 ( .A1(n20967), .A2(n10516), .ZN(n10514) );
INV_X1 U19979 ( .A(n10144), .ZN(n20967) );
NAND2_X1 U19980 ( .A1(n5167), .A2(n5178), .ZN(n5141) );
NAND2_X1 U19981 ( .A1(n10204), .A2(n15816), .ZN(n5583) );
NAND2_X1 U19982 ( .A1(n10068), .A2(n20938), .ZN(n1416) );
NOR2_X1 U19983 ( .A1(n20975), .A2(n10070), .ZN(n10068) );
NAND2_X1 U19984 ( .A1(n20996), .A2(n1580), .ZN(n1501) );
NAND2_X1 U19985 ( .A1(n10541), .A2(n10542), .ZN(n10234) );
AND2_X1 U19986 ( .A1(n15910), .A2(n10230), .ZN(n10542) );
NOR2_X1 U19987 ( .A1(n15912), .A2(n15814), .ZN(n10541) );
NAND2_X1 U19988 ( .A1(n15810), .A2(n15893), .ZN(n10175) );
NOR2_X1 U19989 ( .A1(n20905), .A2(n3042), .ZN(n3590) );
NOR2_X1 U19990 ( .A1(n3566), .A2(n3042), .ZN(n3565) );
NOR2_X1 U19991 ( .A1(n15803), .A2(n19884), .ZN(n3566) );
NAND2_X1 U19992 ( .A1(n2720), .A2(n2591), .ZN(n2655) );
NAND2_X1 U19993 ( .A1(n2723), .A2(n2399), .ZN(n2060) );
NAND2_X1 U19994 ( .A1(n2696), .A2(n2724), .ZN(n2723) );
OR2_X1 U19995 ( .A1(n2440), .A2(n2397), .ZN(n2724) );
NOR2_X1 U19996 ( .A1(n4056), .A2(n5152), .ZN(n5148) );
NOR2_X1 U19997 ( .A1(n16450), .A2(n15806), .ZN(n2271) );
NOR2_X1 U19998 ( .A1(n16450), .A2(n15809), .ZN(n2320) );
NOR2_X1 U19999 ( .A1(n16450), .A2(n15890), .ZN(n2358) );
NAND2_X1 U20000 ( .A1(n16451), .A2(n2727), .ZN(n2448) );
NOR2_X1 U20001 ( .A1(n16450), .A2(n15793), .ZN(n3570) );
NOR2_X1 U20002 ( .A1(n16450), .A2(n15889), .ZN(n2305) );
NOR2_X1 U20003 ( .A1(n16450), .A2(n15885), .ZN(n2259) );
NOR2_X1 U20004 ( .A1(n16450), .A2(n15826), .ZN(n2390) );
NOR2_X1 U20005 ( .A1(n5258), .A2(n1431), .ZN(n5256) );
NOR2_X1 U20006 ( .A1(n4288), .A2(n15906), .ZN(n4933) );
NOR2_X1 U20007 ( .A1(n4288), .A2(n15875), .ZN(n4457) );
NOR2_X1 U20008 ( .A1(n16420), .A2(n15896), .ZN(n4905) );
NOR2_X1 U20009 ( .A1(n4288), .A2(n15897), .ZN(n4886) );
NOR2_X1 U20010 ( .A1(n16420), .A2(n15880), .ZN(n4867) );
NOR2_X1 U20011 ( .A1(n4288), .A2(n15881), .ZN(n4848) );
NOR2_X1 U20012 ( .A1(n16420), .A2(n15882), .ZN(n4829) );
NOR2_X1 U20013 ( .A1(n4288), .A2(n15883), .ZN(n4810) );
NOR2_X1 U20014 ( .A1(n16420), .A2(n15861), .ZN(n4788) );
NOR2_X1 U20015 ( .A1(n4288), .A2(n15862), .ZN(n4767) );
NOR2_X1 U20016 ( .A1(n16420), .A2(n15863), .ZN(n4746) );
NOR2_X1 U20017 ( .A1(n4288), .A2(n15864), .ZN(n4707) );
NOR2_X1 U20018 ( .A1(n4288), .A2(n15865), .ZN(n4686) );
NOR2_X1 U20019 ( .A1(n4288), .A2(n15866), .ZN(n4665) );
NOR2_X1 U20020 ( .A1(n4288), .A2(n15867), .ZN(n4644) );
NOR2_X1 U20021 ( .A1(n4288), .A2(n15868), .ZN(n4623) );
NOR2_X1 U20022 ( .A1(n4288), .A2(n15869), .ZN(n4602) );
NOR2_X1 U20023 ( .A1(n16420), .A2(n15870), .ZN(n4581) );
NOR2_X1 U20024 ( .A1(n4288), .A2(n15871), .ZN(n4560) );
NOR2_X1 U20025 ( .A1(n16420), .A2(n15872), .ZN(n4539) );
NOR2_X1 U20026 ( .A1(n4288), .A2(n15873), .ZN(n4518) );
NOR2_X1 U20027 ( .A1(n16420), .A2(n15874), .ZN(n4478) );
NOR2_X1 U20028 ( .A1(n4288), .A2(n15898), .ZN(n4497) );
NAND2_X1 U20029 ( .A1(n2432), .A2(n2727), .ZN(n2399) );
NAND2_X1 U20030 ( .A1(n10461), .A2(n15798), .ZN(n4051) );
INV_X1 U20031 ( .A(n5237), .ZN(n20923) );
NOR2_X1 U20032 ( .A1(n3579), .A2(n15803), .ZN(n3577) );
NOR2_X1 U20033 ( .A1(n3580), .A2(n3042), .ZN(n3579) );
NOR2_X1 U20034 ( .A1(n3581), .A2(n16457), .ZN(n3580) );
NOR2_X1 U20035 ( .A1(n3582), .A2(n20905), .ZN(n3581) );
NAND2_X1 U20036 ( .A1(n20994), .A2(n10138), .ZN(n10134) );
NAND2_X1 U20037 ( .A1(n10139), .A2(n10140), .ZN(n10138) );
AND2_X1 U20038 ( .A1(n10145), .A2(n10146), .ZN(n10139) );
NOR2_X1 U20039 ( .A1(n10141), .A2(n10142), .ZN(n10140) );
NAND2_X1 U20040 ( .A1(n2814), .A2(n19912), .ZN(n2697) );
NOR2_X1 U20041 ( .A1(n19910), .A2(n2035), .ZN(n2814) );
NOR2_X1 U20042 ( .A1(n2103), .A2(n2518), .ZN(n2517) );
NAND2_X1 U20043 ( .A1(n19906), .A2(n2275), .ZN(n2518) );
AND2_X1 U20044 ( .A1(n7875), .A2(n7722), .ZN(n16262) );
NOR2_X1 U20045 ( .A1(n4960), .A2(n4412), .ZN(n4944) );
NOR2_X1 U20046 ( .A1(n4961), .A2(n4962), .ZN(n4960) );
NAND2_X1 U20047 ( .A1(n4963), .A2(n4964), .ZN(n4962) );
NAND2_X1 U20048 ( .A1(n4975), .A2(n4411), .ZN(n4961) );
NOR2_X1 U20049 ( .A1(n4427), .A2(n4412), .ZN(n4415) );
NOR2_X1 U20050 ( .A1(n4428), .A2(n20918), .ZN(n4427) );
INV_X1 U20051 ( .A(n4411), .ZN(n20918) );
NOR2_X1 U20052 ( .A1(n4430), .A2(n4431), .ZN(n4428) );
NOR2_X1 U20053 ( .A1(n2519), .A2(n2409), .ZN(n2516) );
NOR2_X1 U20054 ( .A1(n20752), .A2(n5385), .ZN(n5427) );
NOR2_X1 U20055 ( .A1(n20214), .A2(n5385), .ZN(n5432) );
NOR2_X1 U20056 ( .A1(n20252), .A2(n16414), .ZN(n5437) );
NOR2_X1 U20057 ( .A1(n20369), .A2(n5385), .ZN(n5450) );
NOR2_X1 U20058 ( .A1(n20608), .A2(n5385), .ZN(n5479) );
NOR2_X1 U20059 ( .A1(n20646), .A2(n5385), .ZN(n5484) );
NOR2_X1 U20060 ( .A1(n20680), .A2(n5385), .ZN(n5489) );
NOR2_X1 U20061 ( .A1(n20687), .A2(n5385), .ZN(n5494) );
NOR2_X1 U20062 ( .A1(n20691), .A2(n5385), .ZN(n5499) );
NOR2_X1 U20063 ( .A1(n20695), .A2(n5385), .ZN(n5504) );
NOR2_X1 U20064 ( .A1(n20707), .A2(n5385), .ZN(n5517) );
NOR2_X1 U20065 ( .A1(n20711), .A2(n16414), .ZN(n5522) );
NOR2_X1 U20066 ( .A1(n20760), .A2(n5385), .ZN(n5527) );
NOR2_X1 U20067 ( .A1(n20865), .A2(n4066), .ZN(n4120) );
NOR2_X1 U20068 ( .A1(n20870), .A2(n4066), .ZN(n4186) );
NOR2_X1 U20069 ( .A1(n20829), .A2(n4066), .ZN(n4240) );
NOR2_X1 U20070 ( .A1(n20831), .A2(n4066), .ZN(n4246) );
NOR2_X1 U20071 ( .A1(n20872), .A2(n4066), .ZN(n4254) );
INV_X1 U20072 ( .A(n1326), .ZN(n21017) );
NOR2_X1 U20073 ( .A1(n1434), .A2(n1435), .ZN(n1433) );
NOR2_X1 U20074 ( .A1(n1436), .A2(n1437), .ZN(n1434) );
NAND2_X1 U20075 ( .A1(n1438), .A2(n1439), .ZN(n1437) );
NOR2_X1 U20076 ( .A1(n1442), .A2(n1443), .ZN(n1436) );
NAND2_X1 U20077 ( .A1(n5578), .A2(n5579), .ZN(n5571) );
NOR2_X1 U20078 ( .A1(n5580), .A2(n5581), .ZN(n5579) );
NOR2_X1 U20079 ( .A1(n5583), .A2(n1431), .ZN(n5578) );
NAND2_X1 U20080 ( .A1(n20963), .A2(n20912), .ZN(n5581) );
INV_X1 U20081 ( .A(n2275), .ZN(n19919) );
NOR2_X1 U20082 ( .A1(n1549), .A2(n1550), .ZN(n1547) );
AND2_X1 U20083 ( .A1(n5127), .A2(n5151), .ZN(n5202) );
NOR2_X1 U20084 ( .A1(n2753), .A2(n3129), .ZN(n3559) );
NOR2_X1 U20085 ( .A1(n2753), .A2(n16434), .ZN(n3573) );
NOR2_X1 U20086 ( .A1(n10185), .A2(n20970), .ZN(n10184) );
NOR2_X1 U20087 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N220), .A2(n5060), .ZN(n5037) );
NOR2_X1 U20088 ( .A1(n5061), .A2(n5062), .ZN(n5060) );
NOR2_X1 U20089 ( .A1(n5063), .A2(n5064), .ZN(n5062) );
NOR2_X1 U20090 ( .A1(n5072), .A2(n5073), .ZN(n5061) );
NOR2_X1 U20091 ( .A1(n8819), .A2(n15890), .ZN(n9963) );
NOR2_X1 U20092 ( .A1(n8819), .A2(n15889), .ZN(n9889) );
NOR2_X1 U20093 ( .A1(n4998), .A2(n16089), .ZN(n4994) );
NOR2_X1 U20094 ( .A1(n4998), .A2(n16086), .ZN(n5022) );
NOR2_X1 U20095 ( .A1(n4998), .A2(n16084), .ZN(n5028) );
NOR2_X1 U20096 ( .A1(n4941), .A2(n5105), .ZN(n5094) );
NAND2_X1 U20097 ( .A1(n4435), .A2(n4940), .ZN(n5105) );
NOR2_X1 U20098 ( .A1(n21009), .A2(n16088), .ZN(n5017) );
NOR2_X1 U20099 ( .A1(n21007), .A2(n16083), .ZN(n5068) );
NOR2_X1 U20100 ( .A1(n21007), .A2(n16091), .ZN(n4988) );
NAND2_X1 U20101 ( .A1(n10230), .A2(n15912), .ZN(n10523) );
NOR2_X1 U20102 ( .A1(n20993), .A2(n1577), .ZN(n1573) );
NOR2_X1 U20103 ( .A1(n1578), .A2(n1549), .ZN(n1577) );
NOR2_X1 U20104 ( .A1(n1525), .A2(n1579), .ZN(n1578) );
NOR2_X1 U20105 ( .A1(n19884), .A2(n3043), .ZN(n3037) );
NAND2_X1 U20106 ( .A1(n16441), .A2(n15812), .ZN(n3043) );
NOR2_X1 U20107 ( .A1(n15859), .A2(n10225), .ZN(n10220) );
NAND2_X1 U20108 ( .A1(n10102), .A2(n15810), .ZN(n10225) );
NOR2_X1 U20109 ( .A1(n3567), .A2(n3568), .ZN(n3563) );
NOR2_X1 U20110 ( .A1(n3042), .A2(n15803), .ZN(n3568) );
NOR2_X1 U20111 ( .A1(n10493), .A2(n15894), .ZN(n10492) );
NOR2_X1 U20112 ( .A1(n3028), .A2(n3710), .ZN(n3713) );
NOR2_X1 U20113 ( .A1(n10103), .A2(n10104), .ZN(n10100) );
NOR2_X1 U20114 ( .A1(n10169), .A2(n10246), .ZN(n10238) );
NOR2_X1 U20115 ( .A1(n5547), .A2(n5548), .ZN(n5546) );
NAND2_X1 U20116 ( .A1(n5549), .A2(n5550), .ZN(n5548) );
NAND2_X1 U20117 ( .A1(n5541), .A2(n21000), .ZN(n5549) );
NOR2_X1 U20118 ( .A1(n10172), .A2(n10173), .ZN(n10171) );
NOR2_X1 U20119 ( .A1(n5101), .A2(n5102), .ZN(n5100) );
NOR2_X1 U20120 ( .A1(n20085), .A2(n20763), .ZN(n5102) );
NOR2_X1 U20121 ( .A1(n4257), .A2(n5104), .ZN(n5101) );
NOR2_X1 U20122 ( .A1(n4996), .A2(n16090), .ZN(n4995) );
NOR2_X1 U20123 ( .A1(n21009), .A2(n16092), .ZN(n4989) );
NOR2_X1 U20124 ( .A1(n10157), .A2(n15826), .ZN(n10480) );
NOR2_X1 U20125 ( .A1(n10157), .A2(n16082), .ZN(n10476) );
NOR2_X1 U20126 ( .A1(n1597), .A2(n1507), .ZN(n1593) );
NOR2_X1 U20127 ( .A1(n2465), .A2(n2466), .ZN(n2464) );
OR2_X1 U20128 ( .A1(n2172), .A2(n19899), .ZN(n2465) );
NAND2_X1 U20129 ( .A1(n19888), .A2(n2468), .ZN(n2466) );
NAND2_X1 U20130 ( .A1(n19904), .A2(n2136), .ZN(n2468) );
NOR2_X1 U20131 ( .A1(n5537), .A2(n5538), .ZN(n5536) );
NAND2_X1 U20132 ( .A1(n5539), .A2(n4941), .ZN(n5538) );
NOR2_X1 U20133 ( .A1(n4431), .A2(n5542), .ZN(n5537) );
NAND2_X1 U20134 ( .A1(n5540), .A2(n5541), .ZN(n5539) );
NOR2_X1 U20135 ( .A1(n2682), .A2(n2683), .ZN(n2681) );
NAND2_X1 U20136 ( .A1(n2684), .A2(n2685), .ZN(n2683) );
NAND2_X1 U20137 ( .A1(n19899), .A2(n2426), .ZN(n2684) );
NAND2_X1 U20138 ( .A1(n2686), .A2(n19914), .ZN(n2685) );
NOR2_X1 U20139 ( .A1(n10413), .A2(n10414), .ZN(n10412) );
NOR2_X1 U20140 ( .A1(n10415), .A2(n10374), .ZN(n10414) );
NOR2_X1 U20141 ( .A1(n15879), .A2(n10446), .ZN(n10413) );
NOR2_X1 U20142 ( .A1(n10416), .A2(n10417), .ZN(n10415) );
NOR2_X1 U20143 ( .A1(n10371), .A2(n1442), .ZN(n10359) );
NOR2_X1 U20144 ( .A1(n10372), .A2(n10373), .ZN(n10371) );
NOR2_X1 U20145 ( .A1(n10367), .A2(n15804), .ZN(n10373) );
NOR2_X1 U20146 ( .A1(n20975), .A2(n15884), .ZN(n10372) );
NOR2_X1 U20147 ( .A1(n10386), .A2(n1439), .ZN(n10378) );
NOR2_X1 U20148 ( .A1(n10389), .A2(n10286), .ZN(n10386) );
NAND2_X1 U20149 ( .A1(n10287), .A2(n10391), .ZN(n10389) );
NAND2_X1 U20150 ( .A1(n10392), .A2(n15892), .ZN(n10391) );
NOR2_X1 U20151 ( .A1(n15913), .A2(n7717), .ZN(n8138) );
NOR2_X1 U20152 ( .A1(n15817), .A2(n7717), .ZN(n8133) );
NOR2_X1 U20153 ( .A1(n10189), .A2(n10173), .ZN(n10178) );
NOR2_X1 U20154 ( .A1(n10095), .A2(n20946), .ZN(n10189) );
AND2_X1 U20155 ( .A1(n16263), .A2(n1541), .ZN(n1695) );
OR2_X1 U20156 ( .A1(n1501), .A2(n1698), .ZN(n16263) );
NOR2_X1 U20157 ( .A1(n1520), .A2(n19965), .ZN(n1574) );
NOR2_X1 U20158 ( .A1(n10097), .A2(n10098), .ZN(n10096) );
NAND2_X1 U20159 ( .A1(n10099), .A2(n20963), .ZN(n10098) );
NOR2_X1 U20160 ( .A1(n5041), .A2(n5042), .ZN(n5039) );
NOR2_X1 U20161 ( .A1(n5043), .A2(n5044), .ZN(n5042) );
NOR2_X1 U20162 ( .A1(n5052), .A2(n5053), .ZN(n5041) );
NAND2_X1 U20163 ( .A1(n5046), .A2(n5047), .ZN(n5043) );
NOR2_X1 U20164 ( .A1(n4932), .A2(n4953), .ZN(n4952) );
NAND2_X1 U20165 ( .A1(n20110), .A2(n15887), .ZN(n4953) );
NOR2_X1 U20166 ( .A1(n3040), .A2(n3041), .ZN(n3039) );
NOR2_X1 U20167 ( .A1(n16442), .A2(n3042), .ZN(n3040) );
NOR2_X1 U20168 ( .A1(n3593), .A2(n1449), .ZN(n3592) );
NOR2_X1 U20169 ( .A1(n19885), .A2(n15793), .ZN(n3593) );
NOR2_X1 U20170 ( .A1(n15813), .A2(n5138), .ZN(n5244) );
NOR2_X1 U20171 ( .A1(n5254), .A2(n5255), .ZN(n5253) );
NAND2_X1 U20172 ( .A1(n5259), .A2(n5260), .ZN(n5254) );
NAND2_X1 U20173 ( .A1(n5256), .A2(n19985), .ZN(n5255) );
NAND2_X1 U20174 ( .A1(n5261), .A2(n5262), .ZN(n5260) );
NOR2_X1 U20175 ( .A1(n15893), .A2(n10168), .ZN(n10167) );
NAND2_X1 U20176 ( .A1(n10169), .A2(n20952), .ZN(n10168) );
AND2_X1 U20177 ( .A1(n2203), .A2(n16264), .ZN(n2199) );
NAND2_X1 U20178 ( .A1(n2036), .A2(n2202), .ZN(n16264) );
NOR2_X1 U20179 ( .A1(n15913), .A2(n7023), .ZN(n7064) );
NOR2_X1 U20180 ( .A1(n15817), .A2(n16399), .ZN(n7056) );
NAND2_X1 U20181 ( .A1(n2675), .A2(n2042), .ZN(n2388) );
INV_X1 U20182 ( .A(n1550), .ZN(n20998) );
OR2_X1 U20183 ( .A1(n16128), .A2(n10253), .ZN(n10193) );
AND2_X1 U20184 ( .A1(n10283), .A2(n10284), .ZN(n5714) );
NOR2_X1 U20185 ( .A1(n1597), .A2(n10288), .ZN(n10283) );
NOR2_X1 U20186 ( .A1(n10285), .A2(n10286), .ZN(n10284) );
OR2_X1 U20187 ( .A1(n15892), .A2(n1439), .ZN(n10288) );
INV_X1 U20188 ( .A(n2308), .ZN(n19921) );
NAND2_X1 U20189 ( .A1(n20922), .A2(n5715), .ZN(n5273) );
NAND2_X1 U20190 ( .A1(n15805), .A2(n15858), .ZN(n5715) );
INV_X1 U20191 ( .A(n2051), .ZN(n19925) );
NOR2_X1 U20192 ( .A1(n10244), .A2(n15859), .ZN(n10521) );
NAND2_X1 U20193 ( .A1(n6306), .A2(n10104), .ZN(n10102) );
INV_X1 U20194 ( .A(n5221), .ZN(n20984) );
NOR2_X1 U20195 ( .A1(n7670), .A2(n3726), .ZN(n7669) );
NOR2_X1 U20196 ( .A1(n7701), .A2(n5147), .ZN(n7670) );
NOR2_X1 U20197 ( .A1(n7630), .A2(n7702), .ZN(n7701) );
NAND2_X1 U20198 ( .A1(n7661), .A2(n20916), .ZN(n7702) );
NOR2_X1 U20199 ( .A1(n7597), .A2(n4028), .ZN(n7596) );
NOR2_X1 U20200 ( .A1(n5147), .A2(n7605), .ZN(n7597) );
NOR2_X1 U20201 ( .A1(n2617), .A2(n2618), .ZN(n2616) );
NOR2_X1 U20202 ( .A1(n2152), .A2(n19925), .ZN(n2618) );
NOR2_X1 U20203 ( .A1(n19940), .A2(n2620), .ZN(n2617) );
NAND2_X1 U20204 ( .A1(n2136), .A2(n2269), .ZN(n2620) );
NOR2_X1 U20205 ( .A1(n5123), .A2(n5124), .ZN(n5122) );
NOR2_X1 U20206 ( .A1(n5126), .A2(n5120), .ZN(n5123) );
NOR2_X1 U20207 ( .A1(n5125), .A2(n4056), .ZN(n5124) );
NOR2_X1 U20208 ( .A1(n5127), .A2(n5128), .ZN(n5126) );
NOR2_X1 U20209 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N220), .A2(n5000), .ZN(n4983) );
NOR2_X1 U20210 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N219), .A2(n5001), .ZN(n5000) );
NOR2_X1 U20211 ( .A1(n5002), .A2(n5003), .ZN(n5001) );
NAND2_X1 U20212 ( .A1(n5004), .A2(n5005), .ZN(n5003) );
NOR2_X1 U20213 ( .A1(n15805), .A2(n15876), .ZN(n10384) );
NAND2_X1 U20214 ( .A1(n3995), .A2(n3996), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N15) );
NAND2_X1 U20215 ( .A1(n3402), .A2(n16442), .ZN(n3996) );
NAND2_X1 U20216 ( .A1(n16440), .A2(n15942), .ZN(n3995) );
NAND2_X1 U20217 ( .A1(n3973), .A2(n3974), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N17) );
NAND2_X1 U20218 ( .A1(n3553), .A2(n16442), .ZN(n3974) );
NAND2_X1 U20219 ( .A1(n16440), .A2(n15944), .ZN(n3973) );
NAND2_X1 U20220 ( .A1(n3950), .A2(n3951), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N19) );
NAND2_X1 U20221 ( .A1(n3543), .A2(n16442), .ZN(n3951) );
NAND2_X1 U20222 ( .A1(n16440), .A2(n15946), .ZN(n3950) );
NAND2_X1 U20223 ( .A1(n3928), .A2(n3929), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N21) );
NAND2_X1 U20224 ( .A1(n3533), .A2(n16442), .ZN(n3929) );
NAND2_X1 U20225 ( .A1(n16440), .A2(n15948), .ZN(n3928) );
NAND2_X1 U20226 ( .A1(n3905), .A2(n3906), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N23) );
NAND2_X1 U20227 ( .A1(n3523), .A2(n16442), .ZN(n3906) );
NAND2_X1 U20228 ( .A1(n16441), .A2(n15950), .ZN(n3905) );
NAND2_X1 U20229 ( .A1(n3883), .A2(n3884), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N25) );
NAND2_X1 U20230 ( .A1(n3513), .A2(n3018), .ZN(n3884) );
NAND2_X1 U20231 ( .A1(n16440), .A2(n15952), .ZN(n3883) );
NAND2_X1 U20232 ( .A1(n3860), .A2(n3861), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N27) );
NAND2_X1 U20233 ( .A1(n3492), .A2(n3018), .ZN(n3861) );
NAND2_X1 U20234 ( .A1(n16440), .A2(n15954), .ZN(n3860) );
NAND2_X1 U20235 ( .A1(n3838), .A2(n3839), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N29) );
NAND2_X1 U20236 ( .A1(n3482), .A2(n3018), .ZN(n3839) );
NAND2_X1 U20237 ( .A1(n16441), .A2(n15956), .ZN(n3838) );
NAND2_X1 U20238 ( .A1(n3816), .A2(n3817), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N31) );
NAND2_X1 U20239 ( .A1(n3472), .A2(n3018), .ZN(n3817) );
NAND2_X1 U20240 ( .A1(n16439), .A2(n15958), .ZN(n3816) );
NAND2_X1 U20241 ( .A1(n3793), .A2(n3794), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N33) );
NAND2_X1 U20242 ( .A1(n3462), .A2(n16442), .ZN(n3794) );
NAND2_X1 U20243 ( .A1(n16440), .A2(n15960), .ZN(n3793) );
NAND2_X1 U20244 ( .A1(n3765), .A2(n3766), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N35) );
NAND2_X1 U20245 ( .A1(n3452), .A2(n16442), .ZN(n3766) );
NAND2_X1 U20246 ( .A1(n16441), .A2(n15962), .ZN(n3765) );
NAND2_X1 U20247 ( .A1(n4032), .A2(n4033), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N11) );
NAND2_X1 U20248 ( .A1(n3422), .A2(n3018), .ZN(n4033) );
NAND2_X1 U20249 ( .A1(n16440), .A2(n15938), .ZN(n4032) );
NAND2_X1 U20250 ( .A1(n4016), .A2(n4017), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N13) );
NAND2_X1 U20251 ( .A1(n3412), .A2(n16442), .ZN(n4017) );
NAND2_X1 U20252 ( .A1(n16440), .A2(n15940), .ZN(n4016) );
NOR2_X1 U20253 ( .A1(n4425), .A2(n4426), .ZN(n4421) );
NAND2_X1 U20254 ( .A1(n3961), .A2(n3962), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N18) );
NAND2_X1 U20255 ( .A1(n3548), .A2(n16442), .ZN(n3962) );
NAND2_X1 U20256 ( .A1(n16440), .A2(n15945), .ZN(n3961) );
NAND2_X1 U20257 ( .A1(n3939), .A2(n3940), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N20) );
NAND2_X1 U20258 ( .A1(n3538), .A2(n3018), .ZN(n3940) );
NAND2_X1 U20259 ( .A1(n16440), .A2(n15947), .ZN(n3939) );
NAND2_X1 U20260 ( .A1(n3917), .A2(n3918), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N22) );
NAND2_X1 U20261 ( .A1(n3528), .A2(n16442), .ZN(n3918) );
NAND2_X1 U20262 ( .A1(n16440), .A2(n15949), .ZN(n3917) );
NAND2_X1 U20263 ( .A1(n3894), .A2(n3895), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N24) );
NAND2_X1 U20264 ( .A1(n3518), .A2(n16442), .ZN(n3895) );
NAND2_X1 U20265 ( .A1(n16440), .A2(n15951), .ZN(n3894) );
NAND2_X1 U20266 ( .A1(n3872), .A2(n3873), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N26) );
NAND2_X1 U20267 ( .A1(n3508), .A2(n3018), .ZN(n3873) );
NAND2_X1 U20268 ( .A1(n16439), .A2(n15953), .ZN(n3872) );
NAND2_X1 U20269 ( .A1(n3849), .A2(n3850), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N28) );
NAND2_X1 U20270 ( .A1(n3487), .A2(n16442), .ZN(n3850) );
NAND2_X1 U20271 ( .A1(n16440), .A2(n15955), .ZN(n3849) );
NAND2_X1 U20272 ( .A1(n3827), .A2(n3828), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N30) );
NAND2_X1 U20273 ( .A1(n3477), .A2(n3018), .ZN(n3828) );
NAND2_X1 U20274 ( .A1(n16441), .A2(n15957), .ZN(n3827) );
NAND2_X1 U20275 ( .A1(n3804), .A2(n3805), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N32) );
NAND2_X1 U20276 ( .A1(n3467), .A2(n16442), .ZN(n3805) );
NAND2_X1 U20277 ( .A1(n16439), .A2(n15959), .ZN(n3804) );
NAND2_X1 U20278 ( .A1(n3781), .A2(n3782), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N34) );
NAND2_X1 U20279 ( .A1(n3457), .A2(n16442), .ZN(n3782) );
NAND2_X1 U20280 ( .A1(n16440), .A2(n15961), .ZN(n3781) );
NAND2_X1 U20281 ( .A1(n3754), .A2(n3755), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N36) );
NAND2_X1 U20282 ( .A1(n3447), .A2(n3018), .ZN(n3755) );
NAND2_X1 U20283 ( .A1(n16441), .A2(n15963), .ZN(n3754) );
NAND2_X1 U20284 ( .A1(n4024), .A2(n4025), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N12) );
NAND2_X1 U20285 ( .A1(n3417), .A2(n3018), .ZN(n4025) );
NAND2_X1 U20286 ( .A1(n16441), .A2(n15939), .ZN(n4024) );
NAND2_X1 U20287 ( .A1(n4009), .A2(n4010), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N14) );
NAND2_X1 U20288 ( .A1(n3407), .A2(n3018), .ZN(n4010) );
NAND2_X1 U20289 ( .A1(n16440), .A2(n15941), .ZN(n4009) );
NAND2_X1 U20290 ( .A1(n3984), .A2(n3985), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N16) );
NAND2_X1 U20291 ( .A1(n3397), .A2(n16442), .ZN(n3985) );
NAND2_X1 U20292 ( .A1(n16440), .A2(n15943), .ZN(n3984) );
NAND2_X1 U20293 ( .A1(n5706), .A2(n5707), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_1) );
NAND2_X1 U20294 ( .A1(n16412), .A2(n15898), .ZN(n5707) );
NAND2_X1 U20295 ( .A1(n5674), .A2(n15862), .ZN(n5706) );
NAND2_X1 U20296 ( .A1(n5694), .A2(n5695), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_2) );
NAND2_X1 U20297 ( .A1(n16411), .A2(n15899), .ZN(n5695) );
NAND2_X1 U20298 ( .A1(n5674), .A2(n15863), .ZN(n5694) );
NAND2_X1 U20299 ( .A1(n5685), .A2(n5686), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_3) );
NAND2_X1 U20300 ( .A1(n16411), .A2(n15900), .ZN(n5686) );
NAND2_X1 U20301 ( .A1(n5674), .A2(n15864), .ZN(n5685) );
NAND2_X1 U20302 ( .A1(n5683), .A2(n5684), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_4) );
NAND2_X1 U20303 ( .A1(n16411), .A2(n15901), .ZN(n5684) );
NAND2_X1 U20304 ( .A1(n5674), .A2(n15865), .ZN(n5683) );
NAND2_X1 U20305 ( .A1(n5681), .A2(n5682), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_5) );
NAND2_X1 U20306 ( .A1(n16411), .A2(n15902), .ZN(n5682) );
NAND2_X1 U20307 ( .A1(n5674), .A2(n15866), .ZN(n5681) );
NAND2_X1 U20308 ( .A1(n5679), .A2(n5680), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_6) );
NAND2_X1 U20309 ( .A1(n16411), .A2(n15903), .ZN(n5680) );
NAND2_X1 U20310 ( .A1(n5674), .A2(n15867), .ZN(n5679) );
NAND2_X1 U20311 ( .A1(n5677), .A2(n5678), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_7) );
NAND2_X1 U20312 ( .A1(n16411), .A2(n15904), .ZN(n5678) );
NAND2_X1 U20313 ( .A1(n5674), .A2(n15868), .ZN(n5677) );
NAND2_X1 U20314 ( .A1(n5675), .A2(n5676), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_8) );
NAND2_X1 U20315 ( .A1(n16411), .A2(n15905), .ZN(n5676) );
NAND2_X1 U20316 ( .A1(n5674), .A2(n15869), .ZN(n5675) );
NAND2_X1 U20317 ( .A1(n5672), .A2(n5673), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_9) );
NAND2_X1 U20318 ( .A1(n16411), .A2(n15906), .ZN(n5673) );
NAND2_X1 U20319 ( .A1(n5674), .A2(n15870), .ZN(n5672) );
NOR2_X1 U20320 ( .A1(n2500), .A2(n2501), .ZN(n2497) );
NOR2_X1 U20321 ( .A1(n2503), .A2(n2504), .ZN(n2500) );
NOR2_X1 U20322 ( .A1(n16446), .A2(n19908), .ZN(n2501) );
NAND2_X1 U20323 ( .A1(n2505), .A2(crash_dump_o_65_), .ZN(n2504) );
NAND2_X1 U20324 ( .A1(n5733), .A2(n5734), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_0) );
NAND2_X1 U20325 ( .A1(n16411), .A2(n15886), .ZN(n5734) );
NAND2_X1 U20326 ( .A1(n5674), .A2(n15861), .ZN(n5733) );
NAND2_X1 U20327 ( .A1(n5731), .A2(n5732), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_10) );
NAND2_X1 U20328 ( .A1(n16412), .A2(n15896), .ZN(n5732) );
NAND2_X1 U20329 ( .A1(n5674), .A2(n15871), .ZN(n5731) );
NAND2_X1 U20330 ( .A1(n5729), .A2(n5730), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_11) );
NAND2_X1 U20331 ( .A1(n16411), .A2(n15897), .ZN(n5730) );
NAND2_X1 U20332 ( .A1(n5674), .A2(n15872), .ZN(n5729) );
NAND2_X1 U20333 ( .A1(n5727), .A2(n5728), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_12) );
NAND2_X1 U20334 ( .A1(n16412), .A2(n15880), .ZN(n5728) );
NAND2_X1 U20335 ( .A1(n5674), .A2(n15873), .ZN(n5727) );
NAND2_X1 U20336 ( .A1(n5725), .A2(n5726), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_13) );
NAND2_X1 U20337 ( .A1(n16411), .A2(n15881), .ZN(n5726) );
NAND2_X1 U20338 ( .A1(n5674), .A2(n15874), .ZN(n5725) );
NAND2_X1 U20339 ( .A1(n5723), .A2(n5724), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_14) );
NAND2_X1 U20340 ( .A1(n16412), .A2(n15882), .ZN(n5724) );
NAND2_X1 U20341 ( .A1(n5674), .A2(n15875), .ZN(n5723) );
NAND2_X1 U20342 ( .A1(n5721), .A2(n5722), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_15) );
NAND2_X1 U20343 ( .A1(n16411), .A2(n15883), .ZN(n5722) );
NAND2_X1 U20344 ( .A1(n5674), .A2(n15891), .ZN(n5721) );
NAND2_X1 U20345 ( .A1(n5719), .A2(n5720), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_16) );
NAND2_X1 U20346 ( .A1(n20992), .A2(n15930), .ZN(n5719) );
NAND2_X1 U20347 ( .A1(n16412), .A2(n15861), .ZN(n5720) );
NAND2_X1 U20348 ( .A1(n5717), .A2(n5718), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_accum_17) );
NAND2_X1 U20349 ( .A1(n20992), .A2(n15931), .ZN(n5717) );
NAND2_X1 U20350 ( .A1(n16411), .A2(n15862), .ZN(n5718) );
NOR2_X1 U20351 ( .A1(n5129), .A2(n5130), .ZN(n5121) );
NOR2_X1 U20352 ( .A1(n5557), .A2(n5547), .ZN(n5554) );
NOR2_X1 U20353 ( .A1(n5541), .A2(n5556), .ZN(n5557) );
NOR2_X1 U20354 ( .A1(n5048), .A2(n5049), .ZN(n5046) );
NOR2_X1 U20355 ( .A1(n21009), .A2(n16094), .ZN(n5049) );
NOR2_X1 U20356 ( .A1(n21007), .A2(n16093), .ZN(n5048) );
NOR2_X1 U20357 ( .A1(n5160), .A2(n5161), .ZN(n5157) );
NOR2_X1 U20358 ( .A1(n20894), .A2(n5162), .ZN(n5161) );
NOR2_X1 U20359 ( .A1(n20914), .A2(n5164), .ZN(n5160) );
NAND2_X1 U20360 ( .A1(n3743), .A2(n3744), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N37) );
NAND2_X1 U20361 ( .A1(n3437), .A2(n16442), .ZN(n3744) );
NAND2_X1 U20362 ( .A1(n16439), .A2(n15964), .ZN(n3743) );
NOR2_X1 U20363 ( .A1(n10502), .A2(n10503), .ZN(n10497) );
NOR2_X1 U20364 ( .A1(n20953), .A2(n15828), .ZN(n10503) );
NOR2_X1 U20365 ( .A1(n10493), .A2(n10506), .ZN(n10502) );
NAND2_X1 U20366 ( .A1(n10501), .A2(n15894), .ZN(n10506) );
NOR2_X1 U20367 ( .A1(n4970), .A2(n15888), .ZN(n4968) );
NOR2_X1 U20368 ( .A1(n4972), .A2(n16114), .ZN(n4970) );
AND2_X1 U20369 ( .A1(n4435), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_0), .ZN(n4972) );
INV_X1 U20370 ( .A(n2432), .ZN(n19942) );
INV_X1 U20371 ( .A(n1571), .ZN(n20995) );
INV_X1 U20372 ( .A(n2591), .ZN(n19923) );
INV_X1 U20373 ( .A(n1554), .ZN(n20997) );
NAND2_X1 U20374 ( .A1(n4425), .A2(n15886), .ZN(n4963) );
INV_X1 U20375 ( .A(n2166), .ZN(n20902) );
NAND2_X1 U20376 ( .A1(n5089), .A2(n4417), .ZN(n4919) );
NOR2_X1 U20377 ( .A1(n5093), .A2(n4939), .ZN(n5089) );
NOR2_X1 U20378 ( .A1(n5094), .A2(n5095), .ZN(n5093) );
NOR2_X1 U20379 ( .A1(n4423), .A2(n5096), .ZN(n5095) );
INV_X1 U20380 ( .A(n10133), .ZN(n20949) );
BUF_X1 U20381 ( .A(n7023), .Z(n16399) );
NAND2_X1 U20382 ( .A1(n2221), .A2(n2222), .ZN(n2220) );
NAND2_X1 U20383 ( .A1(n19875), .A2(n2223), .ZN(n2221) );
NAND2_X1 U20384 ( .A1(n2224), .A2(n2225), .ZN(n2223) );
NOR2_X1 U20385 ( .A1(n2229), .A2(n2230), .ZN(n2224) );
INV_X1 U20386 ( .A(n10104), .ZN(n20946) );
NAND2_X1 U20387 ( .A1(n19874), .A2(n15803), .ZN(n3263) );
INV_X1 U20388 ( .A(n10187), .ZN(n20973) );
INV_X1 U20389 ( .A(n5556), .ZN(n21000) );
NAND2_X1 U20390 ( .A1(n2026), .A2(n2042), .ZN(n2041) );
INV_X1 U20391 ( .A(n1304), .ZN(n21016) );
OR2_X1 U20392 ( .A1(n1431), .A2(n16125), .ZN(n10266) );
AND2_X1 U20393 ( .A1(n10518), .A2(n10519), .ZN(n10145) );
NAND2_X1 U20394 ( .A1(n10520), .A2(n10521), .ZN(n10519) );
NAND2_X1 U20395 ( .A1(n10524), .A2(n1444), .ZN(n10518) );
NOR2_X1 U20396 ( .A1(n10182), .A2(n10246), .ZN(n10520) );
NAND2_X1 U20397 ( .A1(n1444), .A2(n15804), .ZN(n1443) );
AND2_X1 U20398 ( .A1(n20921), .A2(n4957), .ZN(n1422) );
NAND2_X1 U20399 ( .A1(n4958), .A2(n4959), .ZN(n4957) );
NAND2_X1 U20400 ( .A1(n10465), .A2(n5168), .ZN(n5129) );
AND2_X1 U20401 ( .A1(n5162), .A2(n5221), .ZN(n10465) );
NAND2_X1 U20402 ( .A1(n5180), .A2(n20986), .ZN(n5172) );
NOR2_X1 U20403 ( .A1(n20914), .A2(n5182), .ZN(n5180) );
NAND2_X1 U20404 ( .A1(n10287), .A2(n15807), .ZN(n10285) );
INV_X1 U20405 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_N219), .ZN(n21010) );
NAND2_X1 U20406 ( .A1(n5211), .A2(n5212), .ZN(n3586) );
NOR2_X1 U20407 ( .A1(n5222), .A2(n5141), .ZN(n5211) );
NOR2_X1 U20408 ( .A1(n5213), .A2(n5214), .ZN(n5212) );
NAND2_X1 U20409 ( .A1(n5215), .A2(n4056), .ZN(n5214) );
NAND2_X1 U20410 ( .A1(n10215), .A2(n10216), .ZN(n10197) );
OR2_X1 U20411 ( .A1(n10203), .A2(n10173), .ZN(n10216) );
NAND2_X1 U20412 ( .A1(n20980), .A2(n20952), .ZN(n10215) );
NAND2_X1 U20413 ( .A1(n5716), .A2(n5671), .ZN(n5735) );
NAND2_X1 U20414 ( .A1(n5204), .A2(n5205), .ZN(n5159) );
NOR2_X1 U20415 ( .A1(n5208), .A2(n5183), .ZN(n5204) );
NOR2_X1 U20416 ( .A1(n20989), .A2(n20991), .ZN(n5205) );
NOR2_X1 U20417 ( .A1(n3586), .A2(n5162), .ZN(n5208) );
NAND2_X1 U20418 ( .A1(n9838), .A2(n9839), .ZN(n9837) );
NAND2_X1 U20419 ( .A1(n8883), .A2(n15979), .ZN(n9838) );
NAND2_X1 U20420 ( .A1(n19982), .A2(n8310), .ZN(n9839) );
NAND2_X1 U20421 ( .A1(n21002), .A2(n15887), .ZN(n5096) );
NAND2_X1 U20422 ( .A1(n20981), .A2(n10092), .ZN(n6310) );
NAND2_X1 U20423 ( .A1(n10093), .A2(n10094), .ZN(n10092) );
NOR2_X1 U20424 ( .A1(n10100), .A2(n10101), .ZN(n10093) );
NOR2_X1 U20425 ( .A1(n10095), .A2(n10096), .ZN(n10094) );
NAND2_X1 U20426 ( .A1(n21013), .A2(n1359), .ZN(n897) );
NAND2_X1 U20427 ( .A1(n21016), .A2(n1359), .ZN(n898) );
NAND2_X1 U20428 ( .A1(n10269), .A2(n10270), .ZN(n5115) );
NAND2_X1 U20429 ( .A1(n10271), .A2(n20993), .ZN(n10270) );
NAND2_X1 U20430 ( .A1(n6509), .A2(n10272), .ZN(n10269) );
NOR2_X1 U20431 ( .A1(n19988), .A2(n6509), .ZN(n10271) );
NAND2_X1 U20432 ( .A1(n10436), .A2(n10437), .ZN(n5250) );
NOR2_X1 U20433 ( .A1(n10438), .A2(n10433), .ZN(n10436) );
NOR2_X1 U20434 ( .A1(n15815), .A2(rf_raddr_b_o_2_), .ZN(n10437) );
NAND2_X1 U20435 ( .A1(n10450), .A2(n10451), .ZN(n10330) );
NOR2_X1 U20436 ( .A1(n10070), .A2(n1597), .ZN(n10450) );
NOR2_X1 U20437 ( .A1(n5258), .A2(n10374), .ZN(n10451) );
NAND2_X1 U20438 ( .A1(n2332), .A2(n2426), .ZN(n2568) );
NAND2_X1 U20439 ( .A1(n2332), .A2(n2203), .ZN(n2600) );
INV_X1 U20440 ( .A(n2753), .ZN(n19962) );
NAND2_X1 U20441 ( .A1(n5219), .A2(n5162), .ZN(n5210) );
NAND2_X1 U20442 ( .A1(n5220), .A2(n5198), .ZN(n5219) );
NOR2_X1 U20443 ( .A1(n5221), .A2(n15907), .ZN(n5220) );
INV_X1 U20444 ( .A(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fifo_i_add_146_B_1_), .ZN(n19938) );
NAND2_X1 U20445 ( .A1(n10063), .A2(n10064), .ZN(n5267) );
OR2_X1 U20446 ( .A1(n8557), .A2(n9958), .ZN(n10064) );
NAND2_X1 U20447 ( .A1(n9958), .A2(n8557), .ZN(n10063) );
NAND2_X1 U20448 ( .A1(n3047), .A2(n3048), .ZN(n3036) );
NAND2_X1 U20449 ( .A1(n3049), .A2(n16449), .ZN(n3048) );
NAND2_X1 U20450 ( .A1(n16345), .A2(n15793), .ZN(n3047) );
NOR2_X1 U20451 ( .A1(n3050), .A2(n16442), .ZN(n3049) );
NAND2_X1 U20452 ( .A1(n10210), .A2(n20974), .ZN(n10201) );
NOR2_X1 U20453 ( .A1(n10193), .A2(n10185), .ZN(n10210) );
INV_X1 U20454 ( .A(n2035), .ZN(n19907) );
NAND2_X1 U20455 ( .A1(n10282), .A2(n5714), .ZN(n5716) );
NOR2_X1 U20456 ( .A1(n10289), .A2(n10290), .ZN(n10282) );
NOR2_X1 U20457 ( .A1(n15858), .A2(n15805), .ZN(n10289) );
NAND2_X1 U20458 ( .A1(n20991), .A2(n15800), .ZN(n8078) );
NAND2_X1 U20459 ( .A1(n1569), .A2(n1570), .ZN(n1567) );
NOR2_X1 U20460 ( .A1(n1527), .A2(n1572), .ZN(n1569) );
NOR2_X1 U20461 ( .A1(n1553), .A2(n20997), .ZN(n1570) );
NOR2_X1 U20462 ( .A1(n1573), .A2(n1574), .ZN(n1572) );
NAND2_X1 U20463 ( .A1(n3722), .A2(n3723), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N9) );
NAND2_X1 U20464 ( .A1(n3442), .A2(n16442), .ZN(n3723) );
NAND2_X1 U20465 ( .A1(n16440), .A2(n15937), .ZN(n3722) );
NOR2_X1 U20466 ( .A1(n16266), .A2(n16267), .ZN(n16265) );
AND2_X1 U20467 ( .A1(n16441), .A2(n16126), .ZN(n16266) );
AND2_X1 U20468 ( .A1(n3427), .A2(n16442), .ZN(n16267) );
AND2_X1 U20469 ( .A1(n20998), .A2(n1549), .ZN(n1538) );
NAND2_X1 U20470 ( .A1(n1449), .A2(crash_dump_o_65_), .ZN(n2749) );
AND2_X1 U20471 ( .A1(n10524), .A2(n15814), .ZN(n10141) );
AND2_X1 U20472 ( .A1(n2630), .A2(n2631), .ZN(n2624) );
NOR2_X1 U20473 ( .A1(n2632), .A2(n2633), .ZN(n2631) );
NOR2_X1 U20474 ( .A1(n2635), .A2(n2636), .ZN(n2630) );
NOR2_X1 U20475 ( .A1(n19951), .A2(n2166), .ZN(n2632) );
NAND2_X1 U20476 ( .A1(n7580), .A2(n15932), .ZN(n7588) );
NAND2_X1 U20477 ( .A1(n7580), .A2(n15933), .ZN(n7579) );
NAND2_X1 U20478 ( .A1(n5530), .A2(n4425), .ZN(n5386) );
NOR2_X1 U20479 ( .A1(n5374), .A2(n5104), .ZN(n5530) );
NAND2_X1 U20480 ( .A1(n7722), .A2(n8065), .ZN(n7875) );
NAND2_X1 U20481 ( .A1(n19983), .A2(n16384), .ZN(n8065) );
INV_X1 U20482 ( .A(n3290), .ZN(n19874) );
NAND2_X1 U20483 ( .A1(n20988), .A2(n8056), .ZN(n7872) );
AND2_X1 U20484 ( .A1(n10319), .A2(n20968), .ZN(n5125) );
NOR2_X1 U20485 ( .A1(n5249), .A2(n5182), .ZN(n10319) );
NAND2_X1 U20486 ( .A1(n19873), .A2(n15812), .ZN(n3130) );
INV_X1 U20487 ( .A(n10374), .ZN(n20975) );
AND2_X1 U20488 ( .A1(n20984), .A2(n5200), .ZN(n5169) );
NAND2_X1 U20489 ( .A1(n5201), .A2(n5198), .ZN(n5200) );
NOR2_X1 U20490 ( .A1(n5202), .A2(n15907), .ZN(n5201) );
NAND2_X1 U20491 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N219), .A2(n4985), .ZN(n4984) );
NAND2_X1 U20492 ( .A1(n4986), .A2(n4987), .ZN(n4985) );
NOR2_X1 U20493 ( .A1(n4994), .A2(n4995), .ZN(n4986) );
NOR2_X1 U20494 ( .A1(n4988), .A2(n4989), .ZN(n4987) );
NAND2_X1 U20495 ( .A1(n20936), .A2(n9958), .ZN(n5268) );
BUF_X1 U20496 ( .A(n19748), .Z(n16336) );
AND2_X1 U20497 ( .A1(n3715), .A2(n3716), .ZN(n3027) );
NAND2_X1 U20498 ( .A1(n19886), .A2(n15927), .ZN(n3715) );
NAND2_X1 U20499 ( .A1(n3019), .A2(n15878), .ZN(n3716) );
NAND2_X1 U20500 ( .A1(n10133), .A2(n10134), .ZN(n8600) );
NAND2_X1 U20501 ( .A1(n10230), .A2(n15908), .ZN(n10229) );
NOR2_X1 U20502 ( .A1(n3019), .A2(n3024), .ZN(n15750) );
NOR2_X1 U20503 ( .A1(n3025), .A2(n15878), .ZN(n3024) );
AND2_X1 U20504 ( .A1(n2036), .A2(n2491), .ZN(n2068) );
NAND2_X1 U20505 ( .A1(n19875), .A2(n2203), .ZN(n2491) );
OR2_X1 U20506 ( .A1(n1431), .A2(n6509), .ZN(n5112) );
AND2_X1 U20507 ( .A1(n4281), .A2(n4282), .ZN(n4273) );
NOR2_X1 U20508 ( .A1(n4285), .A2(n4286), .ZN(n4281) );
NAND2_X1 U20509 ( .A1(n16353), .A2(n20715), .ZN(n4282) );
NOR2_X1 U20510 ( .A1(data_addr_o_8_), .A2(n4287), .ZN(n4286) );
NAND2_X1 U20511 ( .A1(n19891), .A2(n2440), .ZN(n2718) );
NAND2_X1 U20512 ( .A1(n2025), .A2(n2043), .ZN(n2040) );
NAND2_X1 U20513 ( .A1(n10173), .A2(n10175), .ZN(n10256) );
NAND2_X1 U20514 ( .A1(n10274), .A2(n1596), .ZN(n6545) );
AND2_X1 U20515 ( .A1(n2815), .A2(n2816), .ZN(n2720) );
NOR2_X1 U20516 ( .A1(n2051), .A2(n2275), .ZN(n2816) );
NOR2_X1 U20517 ( .A1(n2103), .A2(n2308), .ZN(n2815) );
AND2_X1 U20518 ( .A1(n7704), .A2(n7705), .ZN(n7661) );
NAND2_X1 U20519 ( .A1(n20913), .A2(n5245), .ZN(n7704) );
INV_X1 U20520 ( .A(n7605), .ZN(n20913) );
NAND2_X1 U20521 ( .A1(n2440), .A2(n2696), .ZN(n2764) );
NAND2_X1 U20522 ( .A1(n1521), .A2(n1522), .ZN(n1511) );
NOR2_X1 U20523 ( .A1(n1527), .A2(n1528), .ZN(n1521) );
NOR2_X1 U20524 ( .A1(n20995), .A2(n1524), .ZN(n1522) );
OR2_X1 U20525 ( .A1(n1525), .A2(n20998), .ZN(n1524) );
NAND2_X1 U20526 ( .A1(n15877), .A2(n4435), .ZN(n4287) );
AND2_X1 U20527 ( .A1(n4400), .A2(n4401), .ZN(n4395) );
NOR2_X1 U20528 ( .A1(n4403), .A2(n4404), .ZN(n4400) );
NAND2_X1 U20529 ( .A1(n16353), .A2(n20746), .ZN(n4401) );
NOR2_X1 U20530 ( .A1(data_addr_o_2_), .A2(n4287), .ZN(n4404) );
AND2_X1 U20531 ( .A1(n4381), .A2(n4382), .ZN(n4376) );
NOR2_X1 U20532 ( .A1(n4384), .A2(n4385), .ZN(n4381) );
NAND2_X1 U20533 ( .A1(n16353), .A2(n20741), .ZN(n4382) );
NOR2_X1 U20534 ( .A1(data_addr_o_3_), .A2(n4287), .ZN(n4385) );
AND2_X1 U20535 ( .A1(n4362), .A2(n4363), .ZN(n4357) );
NOR2_X1 U20536 ( .A1(n4365), .A2(n4366), .ZN(n4362) );
NAND2_X1 U20537 ( .A1(n16353), .A2(n20735), .ZN(n4363) );
NOR2_X1 U20538 ( .A1(data_addr_o_4_), .A2(n16421), .ZN(n4366) );
AND2_X1 U20539 ( .A1(n4343), .A2(n4344), .ZN(n4338) );
NOR2_X1 U20540 ( .A1(n4346), .A2(n4347), .ZN(n4343) );
NAND2_X1 U20541 ( .A1(n16353), .A2(n20730), .ZN(n4344) );
NOR2_X1 U20542 ( .A1(data_addr_o_5_), .A2(n4287), .ZN(n4347) );
AND2_X1 U20543 ( .A1(n4324), .A2(n4325), .ZN(n4319) );
NOR2_X1 U20544 ( .A1(n4327), .A2(n4328), .ZN(n4324) );
NAND2_X1 U20545 ( .A1(n16353), .A2(n20724), .ZN(n4325) );
NOR2_X1 U20546 ( .A1(data_addr_o_6_), .A2(n16421), .ZN(n4328) );
AND2_X1 U20547 ( .A1(n4305), .A2(n4306), .ZN(n4300) );
NOR2_X1 U20548 ( .A1(n4308), .A2(n4309), .ZN(n4305) );
NAND2_X1 U20549 ( .A1(n16353), .A2(n20719), .ZN(n4306) );
NOR2_X1 U20550 ( .A1(data_addr_o_7_), .A2(n4287), .ZN(n4309) );
AND2_X1 U20551 ( .A1(n4929), .A2(n4930), .ZN(n4916) );
NOR2_X1 U20552 ( .A1(n4933), .A2(n4934), .ZN(n4929) );
NAND2_X1 U20553 ( .A1(n20917), .A2(n20711), .ZN(n4930) );
NOR2_X1 U20554 ( .A1(data_addr_o_9_), .A2(n4287), .ZN(n4934) );
AND2_X1 U20555 ( .A1(n4454), .A2(n4455), .ZN(n4449) );
NOR2_X1 U20556 ( .A1(n4457), .A2(n4458), .ZN(n4454) );
NAND2_X1 U20557 ( .A1(n16353), .A2(n20137), .ZN(n4455) );
NOR2_X1 U20558 ( .A1(data_addr_o_30_), .A2(n16421), .ZN(n4458) );
AND2_X1 U20559 ( .A1(n4902), .A2(n4903), .ZN(n4897) );
NOR2_X1 U20560 ( .A1(n4905), .A2(n4906), .ZN(n4902) );
NAND2_X1 U20561 ( .A1(n20917), .A2(n20707), .ZN(n4903) );
NOR2_X1 U20562 ( .A1(data_addr_o_10_), .A2(n4287), .ZN(n4906) );
AND2_X1 U20563 ( .A1(n4883), .A2(n4884), .ZN(n4878) );
NOR2_X1 U20564 ( .A1(n4886), .A2(n4887), .ZN(n4883) );
NAND2_X1 U20565 ( .A1(n20917), .A2(n20703), .ZN(n4884) );
NOR2_X1 U20566 ( .A1(data_addr_o_11_), .A2(n4287), .ZN(n4887) );
AND2_X1 U20567 ( .A1(n4864), .A2(n4865), .ZN(n4859) );
NOR2_X1 U20568 ( .A1(n4867), .A2(n4868), .ZN(n4864) );
NAND2_X1 U20569 ( .A1(n16353), .A2(n20699), .ZN(n4865) );
NOR2_X1 U20570 ( .A1(data_addr_o_12_), .A2(n4287), .ZN(n4868) );
AND2_X1 U20571 ( .A1(n4845), .A2(n4846), .ZN(n4840) );
NOR2_X1 U20572 ( .A1(n4848), .A2(n4849), .ZN(n4845) );
NAND2_X1 U20573 ( .A1(n20917), .A2(n20695), .ZN(n4846) );
NOR2_X1 U20574 ( .A1(data_addr_o_13_), .A2(n4287), .ZN(n4849) );
AND2_X1 U20575 ( .A1(n4826), .A2(n4827), .ZN(n4821) );
NOR2_X1 U20576 ( .A1(n4829), .A2(n4830), .ZN(n4826) );
NAND2_X1 U20577 ( .A1(n16353), .A2(n20691), .ZN(n4827) );
NOR2_X1 U20578 ( .A1(data_addr_o_14_), .A2(n16421), .ZN(n4830) );
AND2_X1 U20579 ( .A1(n4807), .A2(n4808), .ZN(n4802) );
NOR2_X1 U20580 ( .A1(n4810), .A2(n4811), .ZN(n4807) );
NAND2_X1 U20581 ( .A1(n20917), .A2(n20687), .ZN(n4808) );
NOR2_X1 U20582 ( .A1(data_addr_o_15_), .A2(n4287), .ZN(n4811) );
AND2_X1 U20583 ( .A1(n4785), .A2(n4786), .ZN(n4780) );
NOR2_X1 U20584 ( .A1(n4788), .A2(n4789), .ZN(n4785) );
NAND2_X1 U20585 ( .A1(n20917), .A2(n20680), .ZN(n4786) );
NOR2_X1 U20586 ( .A1(data_addr_o_16_), .A2(n4287), .ZN(n4789) );
AND2_X1 U20587 ( .A1(n4764), .A2(n4765), .ZN(n4759) );
NOR2_X1 U20588 ( .A1(n4767), .A2(n4768), .ZN(n4764) );
NAND2_X1 U20589 ( .A1(n20917), .A2(n20646), .ZN(n4765) );
NOR2_X1 U20590 ( .A1(data_addr_o_17_), .A2(n4287), .ZN(n4768) );
AND2_X1 U20591 ( .A1(n4743), .A2(n4744), .ZN(n4738) );
NOR2_X1 U20592 ( .A1(n4746), .A2(n4747), .ZN(n4743) );
NAND2_X1 U20593 ( .A1(n20917), .A2(n20608), .ZN(n4744) );
NOR2_X1 U20594 ( .A1(data_addr_o_18_), .A2(n16421), .ZN(n4747) );
AND2_X1 U20595 ( .A1(n4704), .A2(n4705), .ZN(n4699) );
NOR2_X1 U20596 ( .A1(n4707), .A2(n4708), .ZN(n4704) );
NAND2_X1 U20597 ( .A1(n20917), .A2(n20568), .ZN(n4705) );
NOR2_X1 U20598 ( .A1(data_addr_o_19_), .A2(n4287), .ZN(n4708) );
AND2_X1 U20599 ( .A1(n4683), .A2(n4684), .ZN(n4678) );
NOR2_X1 U20600 ( .A1(n4686), .A2(n4687), .ZN(n4683) );
NAND2_X1 U20601 ( .A1(n20917), .A2(n20528), .ZN(n4684) );
NOR2_X1 U20602 ( .A1(data_addr_o_20_), .A2(n16421), .ZN(n4687) );
AND2_X1 U20603 ( .A1(n4662), .A2(n4663), .ZN(n4657) );
NOR2_X1 U20604 ( .A1(n4665), .A2(n4666), .ZN(n4662) );
NAND2_X1 U20605 ( .A1(n20917), .A2(n20488), .ZN(n4663) );
NOR2_X1 U20606 ( .A1(data_addr_o_21_), .A2(n16421), .ZN(n4666) );
AND2_X1 U20607 ( .A1(n4641), .A2(n4642), .ZN(n4636) );
NOR2_X1 U20608 ( .A1(n4644), .A2(n4645), .ZN(n4641) );
NAND2_X1 U20609 ( .A1(n16353), .A2(n20448), .ZN(n4642) );
NOR2_X1 U20610 ( .A1(data_addr_o_22_), .A2(n16421), .ZN(n4645) );
AND2_X1 U20611 ( .A1(n4620), .A2(n4621), .ZN(n4615) );
NOR2_X1 U20612 ( .A1(n4623), .A2(n4624), .ZN(n4620) );
NAND2_X1 U20613 ( .A1(n20917), .A2(n20408), .ZN(n4621) );
NOR2_X1 U20614 ( .A1(data_addr_o_23_), .A2(n16421), .ZN(n4624) );
AND2_X1 U20615 ( .A1(n4599), .A2(n4600), .ZN(n4594) );
NOR2_X1 U20616 ( .A1(n4602), .A2(n4603), .ZN(n4599) );
NAND2_X1 U20617 ( .A1(n20917), .A2(n20369), .ZN(n4600) );
NOR2_X1 U20618 ( .A1(data_addr_o_24_), .A2(n16421), .ZN(n4603) );
AND2_X1 U20619 ( .A1(n4578), .A2(n4579), .ZN(n4573) );
NOR2_X1 U20620 ( .A1(n4581), .A2(n4582), .ZN(n4578) );
NAND2_X1 U20621 ( .A1(n20917), .A2(n20330), .ZN(n4579) );
NOR2_X1 U20622 ( .A1(data_addr_o_25_), .A2(n16421), .ZN(n4582) );
AND2_X1 U20623 ( .A1(n4557), .A2(n4558), .ZN(n4552) );
NOR2_X1 U20624 ( .A1(n4560), .A2(n4561), .ZN(n4557) );
NAND2_X1 U20625 ( .A1(n16353), .A2(n20291), .ZN(n4558) );
NOR2_X1 U20626 ( .A1(data_addr_o_26_), .A2(n16421), .ZN(n4561) );
AND2_X1 U20627 ( .A1(n4536), .A2(n4537), .ZN(n4531) );
NOR2_X1 U20628 ( .A1(n4539), .A2(n4540), .ZN(n4536) );
NAND2_X1 U20629 ( .A1(n16353), .A2(n20252), .ZN(n4537) );
NOR2_X1 U20630 ( .A1(data_addr_o_27_), .A2(n16421), .ZN(n4540) );
AND2_X1 U20631 ( .A1(n4515), .A2(n4516), .ZN(n4510) );
NOR2_X1 U20632 ( .A1(n4518), .A2(n4519), .ZN(n4515) );
NAND2_X1 U20633 ( .A1(n16353), .A2(n20214), .ZN(n4516) );
NOR2_X1 U20634 ( .A1(data_addr_o_28_), .A2(n16421), .ZN(n4519) );
AND2_X1 U20635 ( .A1(n4475), .A2(n4476), .ZN(n4470) );
NOR2_X1 U20636 ( .A1(n4478), .A2(n4479), .ZN(n4475) );
NAND2_X1 U20637 ( .A1(n16353), .A2(n20176), .ZN(n4476) );
NOR2_X1 U20638 ( .A1(data_addr_o_29_), .A2(n16421), .ZN(n4479) );
AND2_X1 U20639 ( .A1(n4723), .A2(n4724), .ZN(n4718) );
NOR2_X1 U20640 ( .A1(n4726), .A2(n4727), .ZN(n4723) );
NAND2_X1 U20641 ( .A1(n20917), .A2(n20756), .ZN(n4724) );
NOR2_X1 U20642 ( .A1(n16420), .A2(n15886), .ZN(n4726) );
AND2_X1 U20643 ( .A1(n4494), .A2(n4495), .ZN(n4489) );
NOR2_X1 U20644 ( .A1(n4497), .A2(n4498), .ZN(n4494) );
NAND2_X1 U20645 ( .A1(n16353), .A2(n20752), .ZN(n4495) );
NOR2_X1 U20646 ( .A1(alu_adder_result_ex_1), .A2(n16421), .ZN(n4498) );
AND2_X1 U20647 ( .A1(n2642), .A2(n2643), .ZN(n2093) );
NAND2_X1 U20648 ( .A1(n19876), .A2(n2644), .ZN(n2643) );
NOR2_X1 U20649 ( .A1(n2645), .A2(n2646), .ZN(n2642) );
NOR2_X1 U20650 ( .A1(n2647), .A2(n2441), .ZN(n2646) );
AND2_X1 U20651 ( .A1(n2511), .A2(n2512), .ZN(n2074) );
NOR2_X1 U20652 ( .A1(n2508), .A2(n2524), .ZN(n2511) );
NAND2_X1 U20653 ( .A1(n2142), .A2(n2513), .ZN(n2512) );
NOR2_X1 U20654 ( .A1(n2519), .A2(n2471), .ZN(n2524) );
AND2_X1 U20655 ( .A1(n2542), .A2(n2543), .ZN(n2081) );
NAND2_X1 U20656 ( .A1(n2544), .A2(n2275), .ZN(n2543) );
NOR2_X1 U20657 ( .A1(n2508), .A2(n2545), .ZN(n2542) );
NOR2_X1 U20658 ( .A1(n2546), .A2(n2117), .ZN(n2545) );
AND2_X1 U20659 ( .A1(n2560), .A2(n2561), .ZN(n2084) );
NOR2_X1 U20660 ( .A1(n2571), .A2(n2572), .ZN(n2560) );
NOR2_X1 U20661 ( .A1(n2562), .A2(n2563), .ZN(n2561) );
AND2_X1 U20662 ( .A1(n2570), .A2(n19876), .ZN(n2572) );
AND2_X1 U20663 ( .A1(n2586), .A2(n2587), .ZN(n2087) );
NOR2_X1 U20664 ( .A1(n2592), .A2(n2593), .ZN(n2586) );
NOR2_X1 U20665 ( .A1(n2588), .A2(n2589), .ZN(n2587) );
AND2_X1 U20666 ( .A1(n2599), .A2(n19876), .ZN(n2592) );
AND2_X1 U20667 ( .A1(n2678), .A2(n2679), .ZN(n2365) );
NAND2_X1 U20668 ( .A1(n19876), .A2(n2437), .ZN(n2679) );
NOR2_X1 U20669 ( .A1(n2139), .A2(n2680), .ZN(n2678) );
NOR2_X1 U20670 ( .A1(n2681), .A2(n19881), .ZN(n2680) );
NAND2_X1 U20671 ( .A1(n7712), .A2(n20923), .ZN(n7705) );
INV_X1 U20672 ( .A(n1580), .ZN(n19988) );
NAND2_X1 U20673 ( .A1(n2261), .A2(n2275), .ZN(n2274) );
NAND2_X1 U20674 ( .A1(n8418), .A2(n8419), .ZN(n8313) );
NOR2_X1 U20675 ( .A1(n15926), .A2(n8429), .ZN(n8418) );
NOR2_X1 U20676 ( .A1(n1431), .A2(n8420), .ZN(n8419) );
NAND2_X1 U20677 ( .A1(n5242), .A2(n19985), .ZN(n8429) );
NAND2_X1 U20678 ( .A1(n19876), .A2(n2035), .ZN(n2361) );
NAND2_X1 U20679 ( .A1(n2275), .A2(n2393), .ZN(n2392) );
NAND2_X1 U20680 ( .A1(n2394), .A2(n2383), .ZN(n2393) );
NOR2_X1 U20681 ( .A1(n19889), .A2(n2404), .ZN(n2394) );
NOR2_X1 U20682 ( .A1(n2405), .A2(n2058), .ZN(n2404) );
NAND2_X1 U20683 ( .A1(n20962), .A2(n4948), .ZN(n4918) );
NAND2_X1 U20684 ( .A1(n4949), .A2(n4950), .ZN(n4948) );
NAND2_X1 U20685 ( .A1(n21001), .A2(n4423), .ZN(n4950) );
NOR2_X1 U20686 ( .A1(n4426), .A2(n4952), .ZN(n4949) );
NAND2_X1 U20687 ( .A1(n15793), .A2(n15970), .ZN(n3599) );
NAND2_X1 U20688 ( .A1(n20915), .A2(n10323), .ZN(n5146) );
OR2_X1 U20689 ( .A1(n5196), .A2(n15813), .ZN(n10323) );
INV_X1 U20690 ( .A(n5152), .ZN(n20914) );
INV_X1 U20691 ( .A(n5238), .ZN(n20916) );
NAND2_X1 U20692 ( .A1(n10540), .A2(n20965), .ZN(n10143) );
NOR2_X1 U20693 ( .A1(n20990), .A2(n10233), .ZN(n10540) );
NAND2_X1 U20694 ( .A1(n20110), .A2(n15877), .ZN(n4288) );
INV_X1 U20695 ( .A(n10182), .ZN(n20981) );
NAND2_X1 U20696 ( .A1(n3730), .A2(n3731), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_N38) );
NAND2_X1 U20697 ( .A1(n3432), .A2(n16442), .ZN(n3731) );
NAND2_X1 U20698 ( .A1(n16441), .A2(n15965), .ZN(n3730) );
NAND2_X1 U20699 ( .A1(n5086), .A2(n20921), .ZN(n1420) );
AND2_X1 U20700 ( .A1(n5087), .A2(n5088), .ZN(n5086) );
NAND2_X1 U20701 ( .A1(n4937), .A2(n4938), .ZN(n4291) );
NOR2_X1 U20702 ( .A1(n20910), .A2(n4941), .ZN(n4937) );
NOR2_X1 U20703 ( .A1(n4939), .A2(n4940), .ZN(n4938) );
INV_X1 U20704 ( .A(n2863), .ZN(n19943) );
INV_X1 U20705 ( .A(n10097), .ZN(n20974) );
AND2_X1 U20706 ( .A1(n5238), .A2(n7019), .ZN(n6708) );
INV_X1 U20707 ( .A(n10099), .ZN(n20970) );
INV_X1 U20708 ( .A(n1305), .ZN(n21013) );
NAND2_X1 U20709 ( .A1(n10099), .A2(n10263), .ZN(n10262) );
OR2_X1 U20710 ( .A1(n10256), .A2(n20980), .ZN(n10263) );
INV_X1 U20711 ( .A(n4926), .ZN(n21004) );
INV_X1 U20712 ( .A(n10272), .ZN(n20920) );
AND2_X1 U20713 ( .A1(n8117), .A2(n20832), .ZN(n7720) );
NOR2_X1 U20714 ( .A1(n20841), .A2(n1297), .ZN(n8117) );
NAND2_X1 U20715 ( .A1(n2453), .A2(n2018), .ZN(n2601) );
NAND2_X1 U20716 ( .A1(n19889), .A2(n2018), .ZN(n2013) );
NAND2_X1 U20717 ( .A1(n6761), .A2(n6762), .ZN(n6760) );
NAND2_X1 U20718 ( .A1(n20875), .A2(n15804), .ZN(n6761) );
NAND2_X1 U20719 ( .A1(n20876), .A2(crash_dump_o_37_), .ZN(n6762) );
NAND2_X1 U20720 ( .A1(n6783), .A2(n6784), .ZN(n6782) );
NAND2_X1 U20721 ( .A1(n20875), .A2(n15884), .ZN(n6783) );
NAND2_X1 U20722 ( .A1(n20876), .A2(crash_dump_o_35_), .ZN(n6784) );
NAND2_X1 U20723 ( .A1(n6815), .A2(n6816), .ZN(n6814) );
NAND2_X1 U20724 ( .A1(n20875), .A2(n15895), .ZN(n6815) );
NAND2_X1 U20725 ( .A1(n20876), .A2(crash_dump_o_34_), .ZN(n6816) );
NAND2_X1 U20726 ( .A1(n6917), .A2(n6918), .ZN(n6916) );
NAND2_X1 U20727 ( .A1(n20875), .A2(n15820), .ZN(n6917) );
NAND2_X1 U20728 ( .A1(n20876), .A2(crash_dump_o_33_), .ZN(n6918) );
NAND2_X1 U20729 ( .A1(n6993), .A2(n6994), .ZN(n6992) );
NAND2_X1 U20730 ( .A1(n20875), .A2(n15858), .ZN(n6993) );
NAND2_X1 U20731 ( .A1(n20876), .A2(crash_dump_o_44_), .ZN(n6994) );
NAND2_X1 U20732 ( .A1(n7028), .A2(n7029), .ZN(n7027) );
NAND2_X1 U20733 ( .A1(n20875), .A2(n15921), .ZN(n7028) );
NAND2_X1 U20734 ( .A1(n20876), .A2(crash_dump_o_32_), .ZN(n7029) );
NAND2_X1 U20735 ( .A1(n6973), .A2(n6974), .ZN(n6972) );
NAND2_X1 U20736 ( .A1(n20875), .A2(n15805), .ZN(n6973) );
NAND2_X1 U20737 ( .A1(n20876), .A2(crash_dump_o_46_), .ZN(n6974) );
NAND2_X1 U20738 ( .A1(n6983), .A2(n6984), .ZN(n6982) );
NAND2_X1 U20739 ( .A1(n20875), .A2(n15879), .ZN(n6983) );
NAND2_X1 U20740 ( .A1(n20876), .A2(crash_dump_o_45_), .ZN(n6984) );
NAND2_X1 U20741 ( .A1(n6750), .A2(n6751), .ZN(n6749) );
NAND2_X1 U20742 ( .A1(n20875), .A2(n15917), .ZN(n6750) );
NAND2_X1 U20743 ( .A1(n20876), .A2(crash_dump_o_38_), .ZN(n6751) );
NAND2_X1 U20744 ( .A1(n6772), .A2(n6773), .ZN(n6771) );
NAND2_X1 U20745 ( .A1(n20875), .A2(n15876), .ZN(n6772) );
NAND2_X1 U20746 ( .A1(n20876), .A2(crash_dump_o_36_), .ZN(n6773) );
NAND2_X1 U20747 ( .A1(n6822), .A2(n6823), .ZN(n6821) );
NAND2_X1 U20748 ( .A1(id_stage_i_controller_i_N286), .A2(n6708), .ZN(n6822) );
NAND2_X1 U20749 ( .A1(n19974), .A2(n6824), .ZN(n6823) );
NAND2_X1 U20750 ( .A1(n21587), .A2(n21586), .ZN(id_stage_i_controller_i_N286) );
NAND2_X1 U20751 ( .A1(n6894), .A2(n6895), .ZN(n6893) );
NAND2_X1 U20752 ( .A1(id_stage_i_controller_i_N278), .A2(n6708), .ZN(n6894) );
NAND2_X1 U20753 ( .A1(n19974), .A2(n6896), .ZN(n6895) );
NAND2_X1 U20754 ( .A1(n21559), .A2(n21558), .ZN(id_stage_i_controller_i_N278) );
NAND2_X1 U20755 ( .A1(n6840), .A2(n6841), .ZN(n6839) );
NAND2_X1 U20756 ( .A1(id_stage_i_controller_i_N284), .A2(n16403), .ZN(n6840) );
NAND2_X1 U20757 ( .A1(n19974), .A2(n6842), .ZN(n6841) );
NAND2_X1 U20758 ( .A1(n21580), .A2(n21579), .ZN(id_stage_i_controller_i_N284) );
NAND2_X1 U20759 ( .A1(n6849), .A2(n6850), .ZN(n6848) );
NAND2_X1 U20760 ( .A1(id_stage_i_controller_i_N283), .A2(n6708), .ZN(n6849) );
NAND2_X1 U20761 ( .A1(n19974), .A2(n6851), .ZN(n6850) );
NAND2_X1 U20762 ( .A1(n21576), .A2(n21575), .ZN(id_stage_i_controller_i_N283) );
NAND2_X1 U20763 ( .A1(n6858), .A2(n6859), .ZN(n6857) );
NAND2_X1 U20764 ( .A1(id_stage_i_controller_i_N282), .A2(n16403), .ZN(n6858) );
NAND2_X1 U20765 ( .A1(n19974), .A2(n6860), .ZN(n6859) );
NAND2_X1 U20766 ( .A1(n21573), .A2(n21572), .ZN(id_stage_i_controller_i_N282) );
NAND2_X1 U20767 ( .A1(n6867), .A2(n6868), .ZN(n6866) );
NAND2_X1 U20768 ( .A1(id_stage_i_controller_i_N281), .A2(n6708), .ZN(n6867) );
NAND2_X1 U20769 ( .A1(n19974), .A2(n6869), .ZN(n6868) );
NAND2_X1 U20770 ( .A1(n21569), .A2(n21568), .ZN(id_stage_i_controller_i_N281) );
NAND2_X1 U20771 ( .A1(n6876), .A2(n6877), .ZN(n6875) );
NAND2_X1 U20772 ( .A1(id_stage_i_controller_i_N280), .A2(n16403), .ZN(n6876) );
NAND2_X1 U20773 ( .A1(n19974), .A2(n6878), .ZN(n6877) );
NAND2_X1 U20774 ( .A1(n21566), .A2(n21565), .ZN(id_stage_i_controller_i_N280) );
NAND2_X1 U20775 ( .A1(n6885), .A2(n6886), .ZN(n6884) );
NAND2_X1 U20776 ( .A1(id_stage_i_controller_i_N279), .A2(n6708), .ZN(n6885) );
NAND2_X1 U20777 ( .A1(n19974), .A2(n6887), .ZN(n6886) );
NAND2_X1 U20778 ( .A1(n21562), .A2(n21561), .ZN(id_stage_i_controller_i_N279) );
NAND2_X1 U20779 ( .A1(n6903), .A2(n6904), .ZN(n6902) );
NAND2_X1 U20780 ( .A1(id_stage_i_controller_i_N277), .A2(n16403), .ZN(n6903) );
NAND2_X1 U20781 ( .A1(n19974), .A2(n6905), .ZN(n6904) );
NAND2_X1 U20782 ( .A1(n21555), .A2(n21554), .ZN(id_stage_i_controller_i_N277) );
NAND2_X1 U20783 ( .A1(n6923), .A2(n6924), .ZN(n6922) );
NAND2_X1 U20784 ( .A1(id_stage_i_controller_i_N276), .A2(n6708), .ZN(n6923) );
NAND2_X1 U20785 ( .A1(n19974), .A2(n6925), .ZN(n6924) );
NAND2_X1 U20786 ( .A1(n21550), .A2(n21549), .ZN(id_stage_i_controller_i_N276) );
NAND2_X1 U20787 ( .A1(n6932), .A2(n6933), .ZN(n6931) );
NAND2_X1 U20788 ( .A1(id_stage_i_controller_i_N275), .A2(n6708), .ZN(n6932) );
NAND2_X1 U20789 ( .A1(n19974), .A2(n6934), .ZN(n6933) );
NAND2_X1 U20790 ( .A1(n21546), .A2(n21545), .ZN(id_stage_i_controller_i_N275) );
NAND2_X1 U20791 ( .A1(n6950), .A2(n6951), .ZN(n6949) );
NAND2_X1 U20792 ( .A1(id_stage_i_controller_i_N273), .A2(n6708), .ZN(n6950) );
NAND2_X1 U20793 ( .A1(n19974), .A2(n6952), .ZN(n6951) );
NAND2_X1 U20794 ( .A1(n21539), .A2(n21538), .ZN(id_stage_i_controller_i_N273) );
NAND2_X1 U20795 ( .A1(n6941), .A2(n6942), .ZN(n6940) );
NAND2_X1 U20796 ( .A1(id_stage_i_controller_i_N274), .A2(n6708), .ZN(n6941) );
NAND2_X1 U20797 ( .A1(n19974), .A2(n6943), .ZN(n6942) );
NAND2_X1 U20798 ( .A1(n21543), .A2(n21542), .ZN(id_stage_i_controller_i_N274) );
NAND2_X1 U20799 ( .A1(n6831), .A2(n6832), .ZN(n6830) );
NAND2_X1 U20800 ( .A1(id_stage_i_controller_i_N285), .A2(n6708), .ZN(n6831) );
NAND2_X1 U20801 ( .A1(n19974), .A2(n6833), .ZN(n6832) );
NAND2_X1 U20802 ( .A1(n21583), .A2(n21582), .ZN(id_stage_i_controller_i_N285) );
NAND2_X1 U20803 ( .A1(n6801), .A2(n6802), .ZN(n6800) );
NAND2_X1 U20804 ( .A1(id_stage_i_controller_i_N287), .A2(n16403), .ZN(n6801) );
NAND2_X1 U20805 ( .A1(n19974), .A2(n6803), .ZN(n6802) );
NAND2_X1 U20806 ( .A1(n21593), .A2(n21592), .ZN(id_stage_i_controller_i_N287) );
NAND2_X1 U20807 ( .A1(n6789), .A2(n6790), .ZN(n6788) );
NAND2_X1 U20808 ( .A1(id_stage_i_controller_i_N288), .A2(n16403), .ZN(n6789) );
NAND2_X1 U20809 ( .A1(n19974), .A2(n6792), .ZN(n6790) );
NAND2_X1 U20810 ( .A1(n21597), .A2(n21596), .ZN(id_stage_i_controller_i_N288) );
NAND2_X1 U20811 ( .A1(n10352), .A2(n20912), .ZN(n10276) );
NOR2_X1 U20812 ( .A1(n10447), .A2(n1442), .ZN(n10352) );
NOR2_X1 U20813 ( .A1(n15858), .A2(n15804), .ZN(n10447) );
NAND2_X1 U20814 ( .A1(n8421), .A2(n5116), .ZN(n8420) );
NAND2_X1 U20815 ( .A1(n8426), .A2(n20933), .ZN(n8421) );
AND2_X1 U20816 ( .A1(n20962), .A2(n4925), .ZN(n4272) );
NAND2_X1 U20817 ( .A1(n4926), .A2(n4927), .ZN(n4925) );
NAND2_X1 U20818 ( .A1(rf_raddr_b_o_0_), .A2(rf_raddr_b_o_2_), .ZN(n10428) );
NAND2_X1 U20819 ( .A1(n15806), .A2(n15885), .ZN(n10073) );
AND2_X1 U20820 ( .A1(n6301), .A2(n5091), .ZN(n6238) );
NAND2_X1 U20821 ( .A1(n4431), .A2(n4941), .ZN(n6301) );
NAND2_X1 U20822 ( .A1(n7552), .A2(n7553), .ZN(n7551) );
NAND2_X1 U20823 ( .A1(n16396), .A2(n7069), .ZN(n7553) );
NAND2_X1 U20824 ( .A1(n16395), .A2(crash_dump_o_75_), .ZN(n7552) );
NAND2_X1 U20825 ( .A1(n7512), .A2(n7513), .ZN(n7511) );
NAND2_X1 U20826 ( .A1(n16396), .A2(n6952), .ZN(n7513) );
NAND2_X1 U20827 ( .A1(n16395), .A2(crash_dump_o_80_), .ZN(n7512) );
NAND2_X1 U20828 ( .A1(n7520), .A2(n7521), .ZN(n7519) );
NAND2_X1 U20829 ( .A1(n16396), .A2(n7237), .ZN(n7521) );
NAND2_X1 U20830 ( .A1(n16395), .A2(crash_dump_o_79_), .ZN(n7520) );
NAND2_X1 U20831 ( .A1(n7528), .A2(n7529), .ZN(n7527) );
NAND2_X1 U20832 ( .A1(n16396), .A2(n7240), .ZN(n7529) );
NAND2_X1 U20833 ( .A1(n16395), .A2(crash_dump_o_78_), .ZN(n7528) );
NAND2_X1 U20834 ( .A1(n7536), .A2(n7537), .ZN(n7535) );
NAND2_X1 U20835 ( .A1(n16396), .A2(n7243), .ZN(n7537) );
NAND2_X1 U20836 ( .A1(n16395), .A2(crash_dump_o_77_), .ZN(n7536) );
NAND2_X1 U20837 ( .A1(n7544), .A2(n7545), .ZN(n7543) );
NAND2_X1 U20838 ( .A1(n16396), .A2(n7068), .ZN(n7545) );
NAND2_X1 U20839 ( .A1(n16395), .A2(crash_dump_o_76_), .ZN(n7544) );
NAND2_X1 U20840 ( .A1(n7560), .A2(n7561), .ZN(n7559) );
NAND2_X1 U20841 ( .A1(n16396), .A2(n7250), .ZN(n7561) );
NAND2_X1 U20842 ( .A1(n16395), .A2(crash_dump_o_74_), .ZN(n7560) );
NAND2_X1 U20843 ( .A1(n10222), .A2(n10150), .ZN(n10221) );
NAND2_X1 U20844 ( .A1(n10223), .A2(n10103), .ZN(n10222) );
NOR2_X1 U20845 ( .A1(n10182), .A2(n10203), .ZN(n10223) );
NAND2_X1 U20846 ( .A1(n19875), .A2(n2280), .ZN(n2273) );
NAND2_X1 U20847 ( .A1(n2281), .A2(n2282), .ZN(n2280) );
NOR2_X1 U20848 ( .A1(n2286), .A2(n2287), .ZN(n2281) );
NOR2_X1 U20849 ( .A1(n2283), .A2(n2284), .ZN(n2282) );
NAND2_X1 U20850 ( .A1(n7376), .A2(n7377), .ZN(n7375) );
NAND2_X1 U20851 ( .A1(n7318), .A2(n6792), .ZN(n7377) );
NAND2_X1 U20852 ( .A1(n7319), .A2(crash_dump_o_95_), .ZN(n7376) );
NAND2_X1 U20853 ( .A1(n7416), .A2(n7417), .ZN(n7415) );
NAND2_X1 U20854 ( .A1(n7318), .A2(n6842), .ZN(n7417) );
NAND2_X1 U20855 ( .A1(n7319), .A2(crash_dump_o_91_), .ZN(n7416) );
NAND2_X1 U20856 ( .A1(n7424), .A2(n7425), .ZN(n7423) );
NAND2_X1 U20857 ( .A1(n16396), .A2(n6851), .ZN(n7425) );
NAND2_X1 U20858 ( .A1(n16395), .A2(crash_dump_o_90_), .ZN(n7424) );
NAND2_X1 U20859 ( .A1(n7432), .A2(n7433), .ZN(n7431) );
NAND2_X1 U20860 ( .A1(n7318), .A2(n6860), .ZN(n7433) );
NAND2_X1 U20861 ( .A1(n7319), .A2(crash_dump_o_89_), .ZN(n7432) );
NAND2_X1 U20862 ( .A1(n7440), .A2(n7441), .ZN(n7439) );
NAND2_X1 U20863 ( .A1(n16396), .A2(n6869), .ZN(n7441) );
NAND2_X1 U20864 ( .A1(n16395), .A2(crash_dump_o_88_), .ZN(n7440) );
NAND2_X1 U20865 ( .A1(n7448), .A2(n7449), .ZN(n7447) );
NAND2_X1 U20866 ( .A1(n16396), .A2(n6878), .ZN(n7449) );
NAND2_X1 U20867 ( .A1(n16395), .A2(crash_dump_o_87_), .ZN(n7448) );
NAND2_X1 U20868 ( .A1(n7456), .A2(n7457), .ZN(n7455) );
NAND2_X1 U20869 ( .A1(n16396), .A2(n6887), .ZN(n7457) );
NAND2_X1 U20870 ( .A1(n16395), .A2(crash_dump_o_86_), .ZN(n7456) );
NAND2_X1 U20871 ( .A1(n7472), .A2(n7473), .ZN(n7471) );
NAND2_X1 U20872 ( .A1(n16396), .A2(n6905), .ZN(n7473) );
NAND2_X1 U20873 ( .A1(n16395), .A2(crash_dump_o_84_), .ZN(n7472) );
NAND2_X1 U20874 ( .A1(n7488), .A2(n7489), .ZN(n7487) );
NAND2_X1 U20875 ( .A1(n16396), .A2(n6925), .ZN(n7489) );
NAND2_X1 U20876 ( .A1(n16395), .A2(crash_dump_o_83_), .ZN(n7488) );
NAND2_X1 U20877 ( .A1(n7496), .A2(n7497), .ZN(n7495) );
NAND2_X1 U20878 ( .A1(n16396), .A2(n6934), .ZN(n7497) );
NAND2_X1 U20879 ( .A1(n16395), .A2(crash_dump_o_82_), .ZN(n7496) );
NAND2_X1 U20880 ( .A1(n7316), .A2(n7317), .ZN(n7315) );
NAND2_X1 U20881 ( .A1(n7318), .A2(n7179), .ZN(n7317) );
NAND2_X1 U20882 ( .A1(n7319), .A2(crash_dump_o_73_), .ZN(n7316) );
NAND2_X1 U20883 ( .A1(n7328), .A2(n7329), .ZN(n7327) );
NAND2_X1 U20884 ( .A1(n7318), .A2(n7182), .ZN(n7329) );
NAND2_X1 U20885 ( .A1(n7319), .A2(crash_dump_o_72_), .ZN(n7328) );
NAND2_X1 U20886 ( .A1(n7344), .A2(n7345), .ZN(n7343) );
NAND2_X1 U20887 ( .A1(n7318), .A2(n7188), .ZN(n7345) );
NAND2_X1 U20888 ( .A1(n7319), .A2(crash_dump_o_70_), .ZN(n7344) );
NAND2_X1 U20889 ( .A1(n7360), .A2(n7361), .ZN(n7359) );
NAND2_X1 U20890 ( .A1(n7318), .A2(n7194), .ZN(n7361) );
NAND2_X1 U20891 ( .A1(n7319), .A2(crash_dump_o_68_), .ZN(n7360) );
NAND2_X1 U20892 ( .A1(n7336), .A2(n7337), .ZN(n7335) );
NAND2_X1 U20893 ( .A1(n7318), .A2(n7185), .ZN(n7337) );
NAND2_X1 U20894 ( .A1(n7319), .A2(crash_dump_o_71_), .ZN(n7336) );
NAND2_X1 U20895 ( .A1(n7368), .A2(n7369), .ZN(n7367) );
NAND2_X1 U20896 ( .A1(n16396), .A2(n7037), .ZN(n7369) );
NAND2_X1 U20897 ( .A1(n16395), .A2(crash_dump_o_67_), .ZN(n7368) );
NAND2_X1 U20898 ( .A1(n7392), .A2(n7393), .ZN(n7391) );
NAND2_X1 U20899 ( .A1(n7318), .A2(n7203), .ZN(n7393) );
NAND2_X1 U20900 ( .A1(n7319), .A2(crash_dump_o_66_), .ZN(n7392) );
NAND2_X1 U20901 ( .A1(n7504), .A2(n7505), .ZN(n7503) );
NAND2_X1 U20902 ( .A1(n16396), .A2(n6943), .ZN(n7505) );
NAND2_X1 U20903 ( .A1(n16395), .A2(crash_dump_o_81_), .ZN(n7504) );
NAND2_X1 U20904 ( .A1(n7480), .A2(n7481), .ZN(n7479) );
NAND2_X1 U20905 ( .A1(n16396), .A2(n7226), .ZN(n7481) );
NAND2_X1 U20906 ( .A1(n16395), .A2(crash_dump_o_65_), .ZN(n7480) );
NAND2_X1 U20907 ( .A1(n7408), .A2(n7409), .ZN(n7407) );
NAND2_X1 U20908 ( .A1(n16396), .A2(n6833), .ZN(n7409) );
NAND2_X1 U20909 ( .A1(n16395), .A2(crash_dump_o_92_), .ZN(n7408) );
NAND2_X1 U20910 ( .A1(n7400), .A2(n7401), .ZN(n7399) );
NAND2_X1 U20911 ( .A1(n7318), .A2(n6824), .ZN(n7401) );
NAND2_X1 U20912 ( .A1(n7319), .A2(crash_dump_o_93_), .ZN(n7400) );
NAND2_X1 U20913 ( .A1(n7464), .A2(n7465), .ZN(n7463) );
NAND2_X1 U20914 ( .A1(n16396), .A2(n6896), .ZN(n7465) );
NAND2_X1 U20915 ( .A1(n16395), .A2(crash_dump_o_85_), .ZN(n7464) );
NAND2_X1 U20916 ( .A1(n7384), .A2(n7385), .ZN(n7383) );
NAND2_X1 U20917 ( .A1(n16396), .A2(n6803), .ZN(n7385) );
NAND2_X1 U20918 ( .A1(n16395), .A2(crash_dump_o_94_), .ZN(n7384) );
NAND2_X1 U20919 ( .A1(n7352), .A2(n7353), .ZN(n7351) );
NAND2_X1 U20920 ( .A1(n7318), .A2(n7191), .ZN(n7353) );
NAND2_X1 U20921 ( .A1(n7319), .A2(crash_dump_o_69_), .ZN(n7352) );
NAND2_X1 U20922 ( .A1(n19875), .A2(n2159), .ZN(n2157) );
NAND2_X1 U20923 ( .A1(n2160), .A2(n2161), .ZN(n2159) );
NOR2_X1 U20924 ( .A1(n2167), .A2(n2168), .ZN(n2160) );
NOR2_X1 U20925 ( .A1(n2162), .A2(n2163), .ZN(n2161) );
NAND2_X1 U20926 ( .A1(n19875), .A2(n2323), .ZN(n2322) );
NAND2_X1 U20927 ( .A1(n2324), .A2(n2325), .ZN(n2323) );
NOR2_X1 U20928 ( .A1(n2326), .A2(n2327), .ZN(n2325) );
NOR2_X1 U20929 ( .A1(n2329), .A2(n2330), .ZN(n2324) );
NAND2_X1 U20930 ( .A1(n10143), .A2(n10144), .ZN(n10142) );
NAND2_X1 U20931 ( .A1(n1440), .A2(n15876), .ZN(n1438) );
NAND2_X1 U20932 ( .A1(n15889), .A2(n15806), .ZN(n10420) );
NAND2_X1 U20933 ( .A1(n2050), .A2(n2051), .ZN(n2044) );
OR2_X1 U20934 ( .A1(n2030), .A2(n19898), .ZN(n2050) );
NAND2_X1 U20935 ( .A1(n2134), .A2(n19879), .ZN(n2133) );
NAND2_X1 U20936 ( .A1(n2135), .A2(n2136), .ZN(n2134) );
OR2_X1 U20937 ( .A1(n2107), .A2(n19878), .ZN(n2135) );
NAND2_X1 U20938 ( .A1(n2100), .A2(n19879), .ZN(n2099) );
NAND2_X1 U20939 ( .A1(n2102), .A2(n2103), .ZN(n2100) );
NAND2_X1 U20940 ( .A1(n2036), .A2(n2104), .ZN(n2102) );
NAND2_X1 U20941 ( .A1(n7046), .A2(n7047), .ZN(n7045) );
NAND2_X1 U20942 ( .A1(n20929), .A2(n15919), .ZN(n7047) );
NAND2_X1 U20943 ( .A1(n20929), .A2(n16081), .ZN(n7046) );
NAND2_X1 U20944 ( .A1(n10357), .A2(n10358), .ZN(n10356) );
NAND2_X1 U20945 ( .A1(n10290), .A2(n6545), .ZN(n10358) );
NOR2_X1 U20946 ( .A1(n10359), .A2(n10360), .ZN(n10357) );
NOR2_X1 U20947 ( .A1(n10361), .A2(n10362), .ZN(n10360) );
NAND2_X1 U20948 ( .A1(n5193), .A2(n5152), .ZN(n5192) );
NAND2_X1 U20949 ( .A1(n5147), .A2(n5197), .ZN(n5193) );
NAND2_X1 U20950 ( .A1(n20986), .A2(n5173), .ZN(n5197) );
NAND2_X1 U20951 ( .A1(n5142), .A2(n20873), .ZN(n5188) );
NAND2_X1 U20952 ( .A1(n4798), .A2(n4799), .ZN(n4793) );
NAND2_X1 U20953 ( .A1(n4800), .A2(n15861), .ZN(n4799) );
NAND2_X1 U20954 ( .A1(n16350), .A2(data_addr_o_16_), .ZN(n4798) );
NAND2_X1 U20955 ( .A1(n4447), .A2(n4801), .ZN(n4800) );
NAND2_X1 U20956 ( .A1(n4776), .A2(n4777), .ZN(n4772) );
NAND2_X1 U20957 ( .A1(n4778), .A2(n15862), .ZN(n4777) );
NAND2_X1 U20958 ( .A1(n20023), .A2(data_addr_o_17_), .ZN(n4776) );
NAND2_X1 U20959 ( .A1(n4447), .A2(n4779), .ZN(n4778) );
NAND2_X1 U20960 ( .A1(n4755), .A2(n4756), .ZN(n4751) );
NAND2_X1 U20961 ( .A1(n4757), .A2(n15863), .ZN(n4756) );
NAND2_X1 U20962 ( .A1(n16350), .A2(data_addr_o_18_), .ZN(n4755) );
NAND2_X1 U20963 ( .A1(n4447), .A2(n4758), .ZN(n4757) );
NAND2_X1 U20964 ( .A1(n4734), .A2(n4735), .ZN(n4730) );
NAND2_X1 U20965 ( .A1(n4736), .A2(n15864), .ZN(n4735) );
NAND2_X1 U20966 ( .A1(n20023), .A2(data_addr_o_19_), .ZN(n4734) );
NAND2_X1 U20967 ( .A1(n4447), .A2(n4737), .ZN(n4736) );
NAND2_X1 U20968 ( .A1(n4695), .A2(n4696), .ZN(n4691) );
NAND2_X1 U20969 ( .A1(n4697), .A2(n15865), .ZN(n4696) );
NAND2_X1 U20970 ( .A1(n16350), .A2(data_addr_o_20_), .ZN(n4695) );
NAND2_X1 U20971 ( .A1(n4447), .A2(n4698), .ZN(n4697) );
NAND2_X1 U20972 ( .A1(n4674), .A2(n4675), .ZN(n4670) );
NAND2_X1 U20973 ( .A1(n4676), .A2(n15866), .ZN(n4675) );
NAND2_X1 U20974 ( .A1(n20023), .A2(data_addr_o_21_), .ZN(n4674) );
NAND2_X1 U20975 ( .A1(n4447), .A2(n4677), .ZN(n4676) );
NAND2_X1 U20976 ( .A1(n4653), .A2(n4654), .ZN(n4649) );
NAND2_X1 U20977 ( .A1(n4655), .A2(n15867), .ZN(n4654) );
NAND2_X1 U20978 ( .A1(n16350), .A2(data_addr_o_22_), .ZN(n4653) );
NAND2_X1 U20979 ( .A1(n4447), .A2(n4656), .ZN(n4655) );
NAND2_X1 U20980 ( .A1(n4632), .A2(n4633), .ZN(n4628) );
NAND2_X1 U20981 ( .A1(n4634), .A2(n15868), .ZN(n4633) );
NAND2_X1 U20982 ( .A1(n20023), .A2(data_addr_o_23_), .ZN(n4632) );
NAND2_X1 U20983 ( .A1(n4447), .A2(n4635), .ZN(n4634) );
NAND2_X1 U20984 ( .A1(n4611), .A2(n4612), .ZN(n4607) );
NAND2_X1 U20985 ( .A1(n4613), .A2(n15869), .ZN(n4612) );
NAND2_X1 U20986 ( .A1(n16350), .A2(data_addr_o_24_), .ZN(n4611) );
NAND2_X1 U20987 ( .A1(n4447), .A2(n4614), .ZN(n4613) );
NAND2_X1 U20988 ( .A1(n4590), .A2(n4591), .ZN(n4586) );
NAND2_X1 U20989 ( .A1(n4592), .A2(n15870), .ZN(n4591) );
NAND2_X1 U20990 ( .A1(n20023), .A2(data_addr_o_25_), .ZN(n4590) );
NAND2_X1 U20991 ( .A1(n4447), .A2(n4593), .ZN(n4592) );
NAND2_X1 U20992 ( .A1(n4569), .A2(n4570), .ZN(n4565) );
NAND2_X1 U20993 ( .A1(n4571), .A2(n15871), .ZN(n4570) );
NAND2_X1 U20994 ( .A1(n16350), .A2(data_addr_o_26_), .ZN(n4569) );
NAND2_X1 U20995 ( .A1(n4447), .A2(n4572), .ZN(n4571) );
NAND2_X1 U20996 ( .A1(n4548), .A2(n4549), .ZN(n4544) );
NAND2_X1 U20997 ( .A1(n4550), .A2(n15872), .ZN(n4549) );
NAND2_X1 U20998 ( .A1(n20023), .A2(data_addr_o_27_), .ZN(n4548) );
NAND2_X1 U20999 ( .A1(n4447), .A2(n4551), .ZN(n4550) );
NAND2_X1 U21000 ( .A1(n4527), .A2(n4528), .ZN(n4523) );
NAND2_X1 U21001 ( .A1(n4529), .A2(n15873), .ZN(n4528) );
NAND2_X1 U21002 ( .A1(n20023), .A2(data_addr_o_28_), .ZN(n4527) );
NAND2_X1 U21003 ( .A1(n4447), .A2(n4530), .ZN(n4529) );
NAND2_X1 U21004 ( .A1(n4506), .A2(n4507), .ZN(n4502) );
NAND2_X1 U21005 ( .A1(n4508), .A2(n15874), .ZN(n4507) );
NAND2_X1 U21006 ( .A1(n20023), .A2(data_addr_o_29_), .ZN(n4506) );
NAND2_X1 U21007 ( .A1(n4447), .A2(n4509), .ZN(n4508) );
NAND2_X1 U21008 ( .A1(n4466), .A2(n4467), .ZN(n4462) );
NAND2_X1 U21009 ( .A1(n4468), .A2(n15875), .ZN(n4467) );
NAND2_X1 U21010 ( .A1(n20023), .A2(data_addr_o_30_), .ZN(n4466) );
NAND2_X1 U21011 ( .A1(n4447), .A2(n4469), .ZN(n4468) );
NAND2_X1 U21012 ( .A1(n4443), .A2(n4444), .ZN(n4438) );
NAND2_X1 U21013 ( .A1(n4445), .A2(n15891), .ZN(n4444) );
NAND2_X1 U21014 ( .A1(n20023), .A2(data_addr_o_31_), .ZN(n4443) );
NAND2_X1 U21015 ( .A1(n4447), .A2(n4448), .ZN(n4445) );
NAND2_X1 U21016 ( .A1(n1559), .A2(n1560), .ZN(n1558) );
NAND2_X1 U21017 ( .A1(n20993), .A2(n1544), .ZN(n1560) );
NOR2_X1 U21018 ( .A1(n20998), .A2(n1548), .ZN(n1559) );
NAND2_X1 U21019 ( .A1(n4874), .A2(n4875), .ZN(n4873) );
NAND2_X1 U21020 ( .A1(n4876), .A2(n15880), .ZN(n4875) );
NAND2_X1 U21021 ( .A1(n16350), .A2(data_addr_o_12_), .ZN(n4874) );
NAND2_X1 U21022 ( .A1(n4270), .A2(n4877), .ZN(n4876) );
NAND2_X1 U21023 ( .A1(n4855), .A2(n4856), .ZN(n4854) );
NAND2_X1 U21024 ( .A1(n4857), .A2(n15881), .ZN(n4856) );
NAND2_X1 U21025 ( .A1(n16350), .A2(data_addr_o_13_), .ZN(n4855) );
NAND2_X1 U21026 ( .A1(n4270), .A2(n4858), .ZN(n4857) );
NAND2_X1 U21027 ( .A1(n4836), .A2(n4837), .ZN(n4835) );
NAND2_X1 U21028 ( .A1(n4838), .A2(n15882), .ZN(n4837) );
NAND2_X1 U21029 ( .A1(n16350), .A2(data_addr_o_14_), .ZN(n4836) );
NAND2_X1 U21030 ( .A1(n4270), .A2(n4839), .ZN(n4838) );
NAND2_X1 U21031 ( .A1(n4817), .A2(n4818), .ZN(n4816) );
NAND2_X1 U21032 ( .A1(n4819), .A2(n15883), .ZN(n4818) );
NAND2_X1 U21033 ( .A1(n16350), .A2(data_addr_o_15_), .ZN(n4817) );
NAND2_X1 U21034 ( .A1(n4270), .A2(n4820), .ZN(n4819) );
NAND2_X1 U21035 ( .A1(n20955), .A2(rf_raddr_b_o_0_), .ZN(n10510) );
NAND2_X1 U21036 ( .A1(n4912), .A2(n4913), .ZN(n4911) );
NAND2_X1 U21037 ( .A1(n4914), .A2(n15896), .ZN(n4913) );
NAND2_X1 U21038 ( .A1(n16350), .A2(data_addr_o_10_), .ZN(n4912) );
NAND2_X1 U21039 ( .A1(n4270), .A2(n4915), .ZN(n4914) );
NAND2_X1 U21040 ( .A1(n4893), .A2(n4894), .ZN(n4892) );
NAND2_X1 U21041 ( .A1(n4895), .A2(n15897), .ZN(n4894) );
NAND2_X1 U21042 ( .A1(n16350), .A2(data_addr_o_11_), .ZN(n4893) );
NAND2_X1 U21043 ( .A1(n4270), .A2(n4896), .ZN(n4895) );
NAND2_X1 U21044 ( .A1(n4714), .A2(n4715), .ZN(n4713) );
NAND2_X1 U21045 ( .A1(n4716), .A2(n15898), .ZN(n4715) );
NAND2_X1 U21046 ( .A1(n16350), .A2(alu_adder_result_ex_1), .ZN(n4714) );
NAND2_X1 U21047 ( .A1(n4270), .A2(n4717), .ZN(n4716) );
NAND2_X1 U21048 ( .A1(n4485), .A2(n4486), .ZN(n4484) );
NAND2_X1 U21049 ( .A1(n4487), .A2(n15899), .ZN(n4486) );
NAND2_X1 U21050 ( .A1(n20023), .A2(data_addr_o_2_), .ZN(n4485) );
NAND2_X1 U21051 ( .A1(n4270), .A2(n4488), .ZN(n4487) );
NAND2_X1 U21052 ( .A1(n4391), .A2(n4392), .ZN(n4390) );
NAND2_X1 U21053 ( .A1(n4393), .A2(n15900), .ZN(n4392) );
NAND2_X1 U21054 ( .A1(n20023), .A2(data_addr_o_3_), .ZN(n4391) );
NAND2_X1 U21055 ( .A1(n4270), .A2(n4394), .ZN(n4393) );
NAND2_X1 U21056 ( .A1(n4372), .A2(n4373), .ZN(n4371) );
NAND2_X1 U21057 ( .A1(n4374), .A2(n15901), .ZN(n4373) );
NAND2_X1 U21058 ( .A1(n16350), .A2(data_addr_o_4_), .ZN(n4372) );
NAND2_X1 U21059 ( .A1(n4270), .A2(n4375), .ZN(n4374) );
NAND2_X1 U21060 ( .A1(n4353), .A2(n4354), .ZN(n4352) );
NAND2_X1 U21061 ( .A1(n4355), .A2(n15902), .ZN(n4354) );
NAND2_X1 U21062 ( .A1(n20023), .A2(data_addr_o_5_), .ZN(n4353) );
NAND2_X1 U21063 ( .A1(n4270), .A2(n4356), .ZN(n4355) );
NAND2_X1 U21064 ( .A1(n4334), .A2(n4335), .ZN(n4333) );
NAND2_X1 U21065 ( .A1(n4336), .A2(n15903), .ZN(n4335) );
NAND2_X1 U21066 ( .A1(n16350), .A2(data_addr_o_6_), .ZN(n4334) );
NAND2_X1 U21067 ( .A1(n4270), .A2(n4337), .ZN(n4336) );
NAND2_X1 U21068 ( .A1(n4315), .A2(n4316), .ZN(n4314) );
NAND2_X1 U21069 ( .A1(n4317), .A2(n15904), .ZN(n4316) );
NAND2_X1 U21070 ( .A1(n20023), .A2(data_addr_o_7_), .ZN(n4315) );
NAND2_X1 U21071 ( .A1(n4270), .A2(n4318), .ZN(n4317) );
NAND2_X1 U21072 ( .A1(n4296), .A2(n4297), .ZN(n4295) );
NAND2_X1 U21073 ( .A1(n4298), .A2(n15905), .ZN(n4297) );
NAND2_X1 U21074 ( .A1(n16350), .A2(data_addr_o_8_), .ZN(n4296) );
NAND2_X1 U21075 ( .A1(n4270), .A2(n4299), .ZN(n4298) );
NAND2_X1 U21076 ( .A1(n4266), .A2(n4267), .ZN(n4265) );
NAND2_X1 U21077 ( .A1(n4268), .A2(n15906), .ZN(n4267) );
NAND2_X1 U21078 ( .A1(n20023), .A2(data_addr_o_9_), .ZN(n4266) );
NAND2_X1 U21079 ( .A1(n4270), .A2(n4271), .ZN(n4268) );
NAND2_X1 U21080 ( .A1(n10180), .A2(n20951), .ZN(n10179) );
INV_X1 U21081 ( .A(n10166), .ZN(n20951) );
NAND2_X1 U21082 ( .A1(n10183), .A2(n10184), .ZN(n10180) );
NOR2_X1 U21083 ( .A1(n10187), .A2(n10188), .ZN(n10183) );
NAND2_X1 U21084 ( .A1(n4423), .A2(n21002), .ZN(n4422) );
NAND2_X1 U21085 ( .A1(n10482), .A2(rf_raddr_b_o_2_), .ZN(n10487) );
NAND2_X1 U21086 ( .A1(n3018), .A2(n15878), .ZN(n3708) );
INV_X1 U21087 ( .A(n10188), .ZN(n20980) );
NAND2_X1 U21088 ( .A1(n19904), .A2(n2599), .ZN(n2598) );
NAND2_X1 U21089 ( .A1(n16124), .A2(n15821), .ZN(n3605) );
NAND2_X1 U21090 ( .A1(n2043), .A2(n2654), .ZN(n2653) );
OR2_X1 U21091 ( .A1(n2453), .A2(n2332), .ZN(n2654) );
NAND2_X1 U21092 ( .A1(n1516), .A2(n1517), .ZN(n1515) );
OR2_X1 U21093 ( .A1(n20022), .A2(n1518), .ZN(n1517) );
NAND2_X1 U21094 ( .A1(n20996), .A2(n16130), .ZN(n1516) );
OR2_X1 U21095 ( .A1(n10939), .A2(n21577), .ZN(n21574) );
OR2_X1 U21096 ( .A1(n10909), .A2(n21570), .ZN(n21567) );
OR2_X1 U21097 ( .A1(n11495), .A2(n21563), .ZN(n21560) );
OR2_X1 U21098 ( .A1(n10864), .A2(n21556), .ZN(n21553) );
OR2_X1 U21099 ( .A1(n10647), .A2(n21547), .ZN(n21544) );
OR2_X1 U21100 ( .A1(n10817), .A2(n21540), .ZN(n21537) );
OR2_X1 U21101 ( .A1(n10969), .A2(n21584), .ZN(n21581) );
NAND2_X1 U21102 ( .A1(n20996), .A2(n19965), .ZN(n1536) );
NAND2_X1 U21103 ( .A1(n15826), .A2(n16082), .ZN(n10442) );
NAND2_X1 U21104 ( .A1(n4981), .A2(n4982), .ZN(n4980) );
NAND2_X1 U21105 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N220), .A2(n5012), .ZN(n4981) );
NAND2_X1 U21106 ( .A1(n4983), .A2(n4984), .ZN(n4982) );
NAND2_X1 U21107 ( .A1(n5013), .A2(n5014), .ZN(n5012) );
NAND2_X1 U21108 ( .A1(n3025), .A2(n20877), .ZN(n3709) );
NAND2_X1 U21109 ( .A1(n21590), .A2(n21589), .ZN(id_stage_i_controller_i_N259) );
OR2_X1 U21110 ( .A1(n10662), .A2(n21588), .ZN(n21589) );
NAND2_X1 U21111 ( .A1(n21588), .A2(n10662), .ZN(n21590) );
NOR2_X1 U21112 ( .A1(n15928), .A2(n11465), .ZN(n21588) );
AND2_X1 U21113 ( .A1(n5235), .A2(n4056), .ZN(n15563) );
NAND2_X1 U21114 ( .A1(n5236), .A2(n5237), .ZN(n5235) );
NOR2_X1 U21115 ( .A1(n15564), .A2(n5238), .ZN(n5236) );
NAND2_X1 U21116 ( .A1(n4976), .A2(n4977), .ZN(n4975) );
NAND2_X1 U21117 ( .A1(n4978), .A2(n4979), .ZN(n4977) );
NAND2_X1 U21118 ( .A1(n4431), .A2(n5081), .ZN(n4976) );
NAND2_X1 U21119 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N221), .A2(n4980), .ZN(n4979) );
NAND2_X1 U21120 ( .A1(n10482), .A2(rf_raddr_b_o_1_), .ZN(n10498) );
NAND2_X1 U21121 ( .A1(n10423), .A2(n10424), .ZN(n10422) );
NOR2_X1 U21122 ( .A1(n20968), .A2(n8426), .ZN(n10423) );
NOR2_X1 U21123 ( .A1(n10425), .A2(n5251), .ZN(n10424) );
NAND2_X1 U21124 ( .A1(n5015), .A2(n5016), .ZN(n5014) );
NOR2_X1 U21125 ( .A1(n5022), .A2(n5023), .ZN(n5015) );
NOR2_X1 U21126 ( .A1(n5017), .A2(n5018), .ZN(n5016) );
NOR2_X1 U21127 ( .A1(n4996), .A2(n16087), .ZN(n5023) );
INV_X1 U21128 ( .A(n4932), .ZN(n20917) );
NAND2_X1 U21129 ( .A1(n16449), .A2(n15966), .ZN(n2498) );
AND2_X1 U21130 ( .A1(n2018), .A2(n2029), .ZN(n2318) );
NAND2_X1 U21131 ( .A1(n5026), .A2(n5027), .ZN(n5013) );
NOR2_X1 U21132 ( .A1(n5033), .A2(n21010), .ZN(n5026) );
NOR2_X1 U21133 ( .A1(n5028), .A2(n5029), .ZN(n5027) );
NOR2_X1 U21134 ( .A1(n4996), .A2(n16085), .ZN(n5033) );
INV_X1 U21135 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_N220), .ZN(n21011) );
NAND2_X1 U21136 ( .A1(n20904), .A2(n15972), .ZN(n2214) );
NAND2_X1 U21137 ( .A1(n20904), .A2(n15971), .ZN(n2125) );
NAND2_X1 U21138 ( .A1(n16449), .A2(n15967), .ZN(n2527) );
NAND2_X1 U21139 ( .A1(n16449), .A2(n15969), .ZN(n2211) );
NAND2_X1 U21140 ( .A1(n16449), .A2(n15968), .ZN(n2120) );
AND2_X1 U21141 ( .A1(n2308), .A2(n2544), .ZN(n2571) );
AND2_X1 U21142 ( .A1(n1449), .A2(n20904), .ZN(n3591) );
AND2_X1 U21143 ( .A1(n4258), .A2(n4941), .ZN(n5555) );
INV_X1 U21144 ( .A(n5151), .ZN(n20894) );
OR2_X1 U21145 ( .A1(n5268), .A2(n5269), .ZN(n5261) );
AND2_X1 U21146 ( .A1(n5167), .A2(n5168), .ZN(n5166) );
NOR2_X1 U21147 ( .A1(n15911), .A2(n5116), .ZN(n15341) );
NAND2_X1 U21148 ( .A1(n7732), .A2(n7733), .ZN(n14957) );
NAND2_X1 U21149 ( .A1(n7725), .A2(n16005), .ZN(n7732) );
NAND2_X1 U21150 ( .A1(n19976), .A2(n7188), .ZN(n7733) );
INV_X1 U21151 ( .A(n3710), .ZN(n20877) );
AND2_X1 U21152 ( .A1(n7662), .A2(n7025), .ZN(n7660) );
NAND2_X1 U21153 ( .A1(n7160), .A2(n7161), .ZN(n14935) );
NAND2_X1 U21154 ( .A1(n7023), .A2(n15932), .ZN(n7161) );
NAND2_X1 U21155 ( .A1(n16400), .A2(n15977), .ZN(n7160) );
NAND2_X1 U21156 ( .A1(n7156), .A2(n7157), .ZN(n14854) );
NAND2_X1 U21157 ( .A1(n16399), .A2(n15933), .ZN(n7157) );
NAND2_X1 U21158 ( .A1(n16400), .A2(n15978), .ZN(n7156) );
INV_X1 U21159 ( .A(n5178), .ZN(n20987) );
INV_X1 U21160 ( .A(n10274), .ZN(n20976) );
NAND2_X1 U21161 ( .A1(n6562), .A2(n6563), .ZN(n15272) );
NOR2_X1 U21162 ( .A1(n6564), .A2(n6565), .ZN(n6562) );
NAND2_X1 U21163 ( .A1(n19971), .A2(n16040), .ZN(n6563) );
NOR2_X1 U21164 ( .A1(n19749), .A2(n6554), .ZN(n6564) );
NAND2_X1 U21165 ( .A1(n6568), .A2(n6569), .ZN(n15271) );
NOR2_X1 U21166 ( .A1(n6570), .A2(n6571), .ZN(n6568) );
NAND2_X1 U21167 ( .A1(n19971), .A2(n16038), .ZN(n6569) );
NOR2_X1 U21168 ( .A1(n19751), .A2(n6554), .ZN(n6570) );
NAND2_X1 U21169 ( .A1(n6574), .A2(n6575), .ZN(n15270) );
NOR2_X1 U21170 ( .A1(n6576), .A2(n6577), .ZN(n6574) );
NAND2_X1 U21171 ( .A1(n19971), .A2(n16037), .ZN(n6575) );
NOR2_X1 U21172 ( .A1(n19753), .A2(n6554), .ZN(n6576) );
NAND2_X1 U21173 ( .A1(n6622), .A2(n6623), .ZN(n15269) );
NOR2_X1 U21174 ( .A1(n6624), .A2(n6625), .ZN(n6622) );
NAND2_X1 U21175 ( .A1(n19971), .A2(n16032), .ZN(n6623) );
NOR2_X1 U21176 ( .A1(n19769), .A2(n6554), .ZN(n6624) );
NAND2_X1 U21177 ( .A1(n6592), .A2(n6593), .ZN(n15201) );
NOR2_X1 U21178 ( .A1(n6594), .A2(n6595), .ZN(n6592) );
NAND2_X1 U21179 ( .A1(n19971), .A2(n16036), .ZN(n6593) );
NOR2_X1 U21180 ( .A1(n19759), .A2(n6554), .ZN(n6594) );
NAND2_X1 U21181 ( .A1(n6604), .A2(n6605), .ZN(n15171) );
NOR2_X1 U21182 ( .A1(n6606), .A2(n6607), .ZN(n6604) );
NAND2_X1 U21183 ( .A1(n19971), .A2(n16035), .ZN(n6605) );
NOR2_X1 U21184 ( .A1(n19763), .A2(n6554), .ZN(n6606) );
NAND2_X1 U21185 ( .A1(n6610), .A2(n6611), .ZN(n15156) );
NOR2_X1 U21186 ( .A1(n6612), .A2(n6613), .ZN(n6610) );
NAND2_X1 U21187 ( .A1(n19971), .A2(n16034), .ZN(n6611) );
NOR2_X1 U21188 ( .A1(n19765), .A2(n6554), .ZN(n6612) );
NAND2_X1 U21189 ( .A1(n6616), .A2(n6617), .ZN(n15141) );
NOR2_X1 U21190 ( .A1(n6618), .A2(n6619), .ZN(n6616) );
NAND2_X1 U21191 ( .A1(n19971), .A2(n16033), .ZN(n6617) );
NOR2_X1 U21192 ( .A1(n19767), .A2(n6554), .ZN(n6618) );
NAND2_X1 U21193 ( .A1(n6634), .A2(n6635), .ZN(n15111) );
NOR2_X1 U21194 ( .A1(n6636), .A2(n6637), .ZN(n6634) );
NAND2_X1 U21195 ( .A1(n19971), .A2(n16031), .ZN(n6635) );
NOR2_X1 U21196 ( .A1(n19773), .A2(n6554), .ZN(n6636) );
NAND2_X1 U21197 ( .A1(n6640), .A2(n6641), .ZN(n15094) );
NOR2_X1 U21198 ( .A1(n6642), .A2(n6643), .ZN(n6640) );
NAND2_X1 U21199 ( .A1(n19971), .A2(n16030), .ZN(n6641) );
NOR2_X1 U21200 ( .A1(n19775), .A2(n6554), .ZN(n6642) );
NAND2_X1 U21201 ( .A1(n6658), .A2(n6659), .ZN(n15064) );
NOR2_X1 U21202 ( .A1(n6660), .A2(n6661), .ZN(n6658) );
NAND2_X1 U21203 ( .A1(n19971), .A2(n16028), .ZN(n6659) );
NOR2_X1 U21204 ( .A1(n19781), .A2(n6554), .ZN(n6660) );
NAND2_X1 U21205 ( .A1(n6664), .A2(n6665), .ZN(n15050) );
NOR2_X1 U21206 ( .A1(n6666), .A2(n6667), .ZN(n6664) );
NAND2_X1 U21207 ( .A1(n19971), .A2(n16027), .ZN(n6665) );
NOR2_X1 U21208 ( .A1(n19783), .A2(n6554), .ZN(n6666) );
NAND2_X1 U21209 ( .A1(n6670), .A2(n6671), .ZN(n15035) );
NOR2_X1 U21210 ( .A1(n6672), .A2(n6673), .ZN(n6670) );
NAND2_X1 U21211 ( .A1(n19971), .A2(n16026), .ZN(n6671) );
NOR2_X1 U21212 ( .A1(n19785), .A2(n6554), .ZN(n6672) );
NAND2_X1 U21213 ( .A1(n6676), .A2(n6677), .ZN(n15019) );
NOR2_X1 U21214 ( .A1(n6678), .A2(n6679), .ZN(n6676) );
NAND2_X1 U21215 ( .A1(n19971), .A2(n16025), .ZN(n6677) );
NOR2_X1 U21216 ( .A1(n19787), .A2(n6554), .ZN(n6678) );
NAND2_X1 U21217 ( .A1(n6688), .A2(n6689), .ZN(n14995) );
NOR2_X1 U21218 ( .A1(n6690), .A2(n6691), .ZN(n6688) );
NAND2_X1 U21219 ( .A1(n19971), .A2(n16024), .ZN(n6689) );
NOR2_X1 U21220 ( .A1(n19791), .A2(n6554), .ZN(n6690) );
NAND2_X1 U21221 ( .A1(n6546), .A2(n6547), .ZN(n14981) );
NOR2_X1 U21222 ( .A1(n6549), .A2(n6550), .ZN(n6546) );
NAND2_X1 U21223 ( .A1(n19971), .A2(n16039), .ZN(n6547) );
NOR2_X1 U21224 ( .A1(n19793), .A2(n6554), .ZN(n6549) );
NAND2_X1 U21225 ( .A1(n6555), .A2(n6556), .ZN(n14967) );
NOR2_X1 U21226 ( .A1(n6557), .A2(n6558), .ZN(n6555) );
NAND2_X1 U21227 ( .A1(n19971), .A2(n16023), .ZN(n6556) );
NOR2_X1 U21228 ( .A1(n19795), .A2(n6554), .ZN(n6557) );
NAND2_X1 U21229 ( .A1(n6646), .A2(n6647), .ZN(n14898) );
NOR2_X1 U21230 ( .A1(n6648), .A2(n6649), .ZN(n6646) );
NAND2_X1 U21231 ( .A1(n19971), .A2(n16029), .ZN(n6647) );
NOR2_X1 U21232 ( .A1(n19777), .A2(n6554), .ZN(n6648) );
NAND2_X1 U21233 ( .A1(n7298), .A2(n7299), .ZN(n15765) );
NAND2_X1 U21234 ( .A1(n19973), .A2(n6833), .ZN(n7298) );
NAND2_X1 U21235 ( .A1(n7257), .A2(n16014), .ZN(n7299) );
NAND2_X1 U21236 ( .A1(n7281), .A2(n7282), .ZN(n15760) );
NAND2_X1 U21237 ( .A1(n19973), .A2(n6943), .ZN(n7281) );
NAND2_X1 U21238 ( .A1(n7257), .A2(n16129), .ZN(n7282) );
NAND2_X1 U21239 ( .A1(n7269), .A2(n7270), .ZN(n15401) );
NAND2_X1 U21240 ( .A1(n19973), .A2(n6896), .ZN(n7269) );
NAND2_X1 U21241 ( .A1(n7257), .A2(n16011), .ZN(n7270) );
NAND2_X1 U21242 ( .A1(n7295), .A2(n7296), .ZN(n15400) );
NAND2_X1 U21243 ( .A1(n19973), .A2(n6824), .ZN(n7295) );
NAND2_X1 U21244 ( .A1(n7257), .A2(n16008), .ZN(n7296) );
NAND2_X1 U21245 ( .A1(n7292), .A2(n7293), .ZN(n15399) );
NAND2_X1 U21246 ( .A1(n19973), .A2(n6803), .ZN(n7292) );
NAND2_X1 U21247 ( .A1(n7257), .A2(n16127), .ZN(n7293) );
NAND2_X1 U21248 ( .A1(n7289), .A2(n7290), .ZN(n15398) );
NAND2_X1 U21249 ( .A1(n19973), .A2(n7069), .ZN(n7289) );
NAND2_X1 U21250 ( .A1(n7257), .A2(n16016), .ZN(n7290) );
NAND2_X1 U21251 ( .A1(n7284), .A2(n7285), .ZN(n15397) );
NAND2_X1 U21252 ( .A1(n19973), .A2(n7037), .ZN(n7284) );
NAND2_X1 U21253 ( .A1(n7257), .A2(n16015), .ZN(n7285) );
NAND2_X1 U21254 ( .A1(n7301), .A2(n7302), .ZN(n15221) );
NAND2_X1 U21255 ( .A1(n19973), .A2(n6842), .ZN(n7301) );
NAND2_X1 U21256 ( .A1(n7257), .A2(n16004), .ZN(n7302) );
NAND2_X1 U21257 ( .A1(n7304), .A2(n7305), .ZN(n15206) );
NAND2_X1 U21258 ( .A1(n19973), .A2(n6851), .ZN(n7304) );
NAND2_X1 U21259 ( .A1(n7257), .A2(n16001), .ZN(n7305) );
NAND2_X1 U21260 ( .A1(n7255), .A2(n7256), .ZN(n15191) );
NAND2_X1 U21261 ( .A1(n19973), .A2(n6860), .ZN(n7255) );
NAND2_X1 U21262 ( .A1(n7257), .A2(n16000), .ZN(n7256) );
NAND2_X1 U21263 ( .A1(n7260), .A2(n7261), .ZN(n15176) );
NAND2_X1 U21264 ( .A1(n19973), .A2(n6869), .ZN(n7260) );
NAND2_X1 U21265 ( .A1(n7257), .A2(n16009), .ZN(n7261) );
NAND2_X1 U21266 ( .A1(n7263), .A2(n7264), .ZN(n15161) );
NAND2_X1 U21267 ( .A1(n19973), .A2(n6878), .ZN(n7263) );
NAND2_X1 U21268 ( .A1(n7257), .A2(n16010), .ZN(n7264) );
NAND2_X1 U21269 ( .A1(n7266), .A2(n7267), .ZN(n15146) );
NAND2_X1 U21270 ( .A1(n19973), .A2(n6887), .ZN(n7266) );
NAND2_X1 U21271 ( .A1(n7257), .A2(n16003), .ZN(n7267) );
NAND2_X1 U21272 ( .A1(n7272), .A2(n7273), .ZN(n15131) );
NAND2_X1 U21273 ( .A1(n19973), .A2(n6905), .ZN(n7272) );
NAND2_X1 U21274 ( .A1(n7257), .A2(n16013), .ZN(n7273) );
NAND2_X1 U21275 ( .A1(n7275), .A2(n7276), .ZN(n15116) );
NAND2_X1 U21276 ( .A1(n19973), .A2(n6925), .ZN(n7275) );
NAND2_X1 U21277 ( .A1(n7257), .A2(n16012), .ZN(n7276) );
NAND2_X1 U21278 ( .A1(n7278), .A2(n7279), .ZN(n15101) );
NAND2_X1 U21279 ( .A1(n19973), .A2(n6934), .ZN(n7278) );
NAND2_X1 U21280 ( .A1(n7257), .A2(n16006), .ZN(n7279) );
NAND2_X1 U21281 ( .A1(n7307), .A2(n7308), .ZN(n15084) );
NAND2_X1 U21282 ( .A1(n19973), .A2(n6952), .ZN(n7307) );
NAND2_X1 U21283 ( .A1(n7257), .A2(n16017), .ZN(n7308) );
NAND2_X1 U21284 ( .A1(n21449), .A2(n21448), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_2) );
OR2_X1 U21285 ( .A1(n21447), .A2(n21446), .ZN(n21449) );
NAND2_X1 U21286 ( .A1(n21447), .A2(n21446), .ZN(n21448) );
AND2_X1 U21287 ( .A1(n21445), .A2(n21444), .ZN(n21447) );
NAND2_X1 U21288 ( .A1(n7777), .A2(n7778), .ZN(n15067) );
NAND2_X1 U21289 ( .A1(n7725), .A2(n16018), .ZN(n7778) );
NAND2_X1 U21290 ( .A1(n19976), .A2(n7237), .ZN(n7777) );
NAND2_X1 U21291 ( .A1(n7780), .A2(n7781), .ZN(n15052) );
NAND2_X1 U21292 ( .A1(n7725), .A2(n16019), .ZN(n7781) );
NAND2_X1 U21293 ( .A1(n19976), .A2(n7240), .ZN(n7780) );
NAND2_X1 U21294 ( .A1(n7783), .A2(n7784), .ZN(n15038) );
NAND2_X1 U21295 ( .A1(n7725), .A2(n16020), .ZN(n7784) );
NAND2_X1 U21296 ( .A1(n16347), .A2(n7243), .ZN(n7783) );
NAND2_X1 U21297 ( .A1(n7790), .A2(n7791), .ZN(n14999) );
NAND2_X1 U21298 ( .A1(n7725), .A2(n16021), .ZN(n7791) );
NAND2_X1 U21299 ( .A1(n19976), .A2(n7250), .ZN(n7790) );
NAND2_X1 U21300 ( .A1(n7723), .A2(n7724), .ZN(n14985) );
NAND2_X1 U21301 ( .A1(n7725), .A2(n16022), .ZN(n7724) );
NAND2_X1 U21302 ( .A1(n19976), .A2(n7179), .ZN(n7723) );
INV_X1 U21303 ( .A(n10433), .ZN(n20969) );
NAND2_X1 U21304 ( .A1(n5551), .A2(n5552), .ZN(n15545) );
NAND2_X1 U21305 ( .A1(n5374), .A2(n15888), .ZN(n5551) );
NAND2_X1 U21306 ( .A1(n20906), .A2(n5553), .ZN(n5552) );
NAND2_X1 U21307 ( .A1(n5554), .A2(n5555), .ZN(n5553) );
INV_X1 U21308 ( .A(n10244), .ZN(n20978) );
NAND2_X1 U21309 ( .A1(n5380), .A2(n5381), .ZN(n15543) );
NOR2_X1 U21310 ( .A1(n5383), .A2(n5384), .ZN(n5380) );
NAND2_X1 U21311 ( .A1(n16415), .A2(n16121), .ZN(n5381) );
NOR2_X1 U21312 ( .A1(n20715), .A2(n16414), .ZN(n5384) );
NAND2_X1 U21313 ( .A1(n5387), .A2(n5388), .ZN(n15542) );
NOR2_X1 U21314 ( .A1(n5390), .A2(n5391), .ZN(n5387) );
NAND2_X1 U21315 ( .A1(n16415), .A2(n16134), .ZN(n5388) );
NOR2_X1 U21316 ( .A1(n20719), .A2(n16414), .ZN(n5391) );
NAND2_X1 U21317 ( .A1(n5392), .A2(n5393), .ZN(n15541) );
NOR2_X1 U21318 ( .A1(n5395), .A2(n5396), .ZN(n5392) );
NAND2_X1 U21319 ( .A1(n16415), .A2(n16135), .ZN(n5393) );
NOR2_X1 U21320 ( .A1(n20724), .A2(n16414), .ZN(n5396) );
NAND2_X1 U21321 ( .A1(n5397), .A2(n5398), .ZN(n15540) );
NOR2_X1 U21322 ( .A1(n5400), .A2(n5401), .ZN(n5397) );
NAND2_X1 U21323 ( .A1(n16415), .A2(n16136), .ZN(n5398) );
NOR2_X1 U21324 ( .A1(n20730), .A2(n16414), .ZN(n5401) );
NAND2_X1 U21325 ( .A1(n5402), .A2(n5403), .ZN(n15539) );
NOR2_X1 U21326 ( .A1(n5404), .A2(n5405), .ZN(n5402) );
NAND2_X1 U21327 ( .A1(n16415), .A2(n16083), .ZN(n5403) );
NOR2_X1 U21328 ( .A1(n20735), .A2(n16414), .ZN(n5405) );
NAND2_X1 U21329 ( .A1(n5406), .A2(n5407), .ZN(n15538) );
NOR2_X1 U21330 ( .A1(n5408), .A2(n5409), .ZN(n5406) );
NAND2_X1 U21331 ( .A1(n16415), .A2(n16122), .ZN(n5407) );
NOR2_X1 U21332 ( .A1(n20741), .A2(n16414), .ZN(n5409) );
NAND2_X1 U21333 ( .A1(n5410), .A2(n5411), .ZN(n15537) );
NOR2_X1 U21334 ( .A1(n5413), .A2(n5414), .ZN(n5410) );
NAND2_X1 U21335 ( .A1(n16415), .A2(n16137), .ZN(n5411) );
NOR2_X1 U21336 ( .A1(n20746), .A2(n16414), .ZN(n5414) );
NAND2_X1 U21337 ( .A1(n5415), .A2(n5416), .ZN(n15536) );
NOR2_X1 U21338 ( .A1(n5417), .A2(n5418), .ZN(n5415) );
NAND2_X1 U21339 ( .A1(n16415), .A2(n16084), .ZN(n5416) );
NOR2_X1 U21340 ( .A1(n20137), .A2(n16414), .ZN(n5418) );
NAND2_X1 U21341 ( .A1(n4059), .A2(n4060), .ZN(n15505) );
NOR2_X1 U21342 ( .A1(n4063), .A2(n4064), .ZN(n4059) );
NAND2_X1 U21343 ( .A1(n4061), .A2(n16138), .ZN(n4060) );
NOR2_X1 U21344 ( .A1(n20834), .A2(n16426), .ZN(n4064) );
NAND2_X1 U21345 ( .A1(n4068), .A2(n4069), .ZN(n15504) );
NOR2_X1 U21346 ( .A1(n4071), .A2(n4072), .ZN(n4068) );
NAND2_X1 U21347 ( .A1(n4061), .A2(n16139), .ZN(n4069) );
NOR2_X1 U21348 ( .A1(n20836), .A2(n16426), .ZN(n4072) );
NAND2_X1 U21349 ( .A1(n4074), .A2(n4075), .ZN(n15503) );
NOR2_X1 U21350 ( .A1(n4077), .A2(n4078), .ZN(n4074) );
NAND2_X1 U21351 ( .A1(n4061), .A2(n16140), .ZN(n4075) );
NOR2_X1 U21352 ( .A1(n20840), .A2(n16426), .ZN(n4078) );
NAND2_X1 U21353 ( .A1(n4080), .A2(n4081), .ZN(n15502) );
NOR2_X1 U21354 ( .A1(n4083), .A2(n4084), .ZN(n4080) );
NAND2_X1 U21355 ( .A1(n16427), .A2(n16141), .ZN(n4081) );
NOR2_X1 U21356 ( .A1(n20842), .A2(n16426), .ZN(n4084) );
NAND2_X1 U21357 ( .A1(n4086), .A2(n4087), .ZN(n15501) );
NOR2_X1 U21358 ( .A1(n4089), .A2(n4090), .ZN(n4086) );
NAND2_X1 U21359 ( .A1(n4061), .A2(n16142), .ZN(n4087) );
NOR2_X1 U21360 ( .A1(n20847), .A2(n16426), .ZN(n4090) );
NAND2_X1 U21361 ( .A1(n4092), .A2(n4093), .ZN(n15500) );
NOR2_X1 U21362 ( .A1(n4095), .A2(n4096), .ZN(n4092) );
NAND2_X1 U21363 ( .A1(n16427), .A2(n16143), .ZN(n4093) );
NOR2_X1 U21364 ( .A1(n20854), .A2(n16426), .ZN(n4096) );
NAND2_X1 U21365 ( .A1(n4098), .A2(n4099), .ZN(n15499) );
NOR2_X1 U21366 ( .A1(n4101), .A2(n4102), .ZN(n4098) );
NAND2_X1 U21367 ( .A1(n4061), .A2(n16144), .ZN(n4099) );
NOR2_X1 U21368 ( .A1(n20862), .A2(n16426), .ZN(n4102) );
NAND2_X1 U21369 ( .A1(n4104), .A2(n4105), .ZN(n15498) );
NOR2_X1 U21370 ( .A1(n4107), .A2(n4108), .ZN(n4104) );
NAND2_X1 U21371 ( .A1(n16427), .A2(n16041), .ZN(n4105) );
NOR2_X1 U21372 ( .A1(n20764), .A2(n16426), .ZN(n4108) );
NAND2_X1 U21373 ( .A1(n3014), .A2(n3015), .ZN(n14834) );
NOR2_X1 U21374 ( .A1(n3016), .A2(n3017), .ZN(n3014) );
NAND2_X1 U21375 ( .A1(n16445), .A2(n15996), .ZN(n3015) );
NOR2_X1 U21376 ( .A1(n19866), .A2(n2901), .ZN(n3016) );
NAND2_X1 U21377 ( .A1(n3006), .A2(n3007), .ZN(n14830) );
NOR2_X1 U21378 ( .A1(n3008), .A2(n3009), .ZN(n3006) );
NAND2_X1 U21379 ( .A1(n16445), .A2(n15991), .ZN(n3007) );
NOR2_X1 U21380 ( .A1(n19861), .A2(n16443), .ZN(n3008) );
NAND2_X1 U21381 ( .A1(n3002), .A2(n3003), .ZN(n14828) );
NOR2_X1 U21382 ( .A1(n3004), .A2(n3005), .ZN(n3002) );
NAND2_X1 U21383 ( .A1(n16445), .A2(n15992), .ZN(n3003) );
NOR2_X1 U21384 ( .A1(n19858), .A2(n2901), .ZN(n3004) );
NAND2_X1 U21385 ( .A1(n2998), .A2(n2999), .ZN(n14826) );
NOR2_X1 U21386 ( .A1(n3000), .A2(n3001), .ZN(n2998) );
NAND2_X1 U21387 ( .A1(n16445), .A2(n15993), .ZN(n2999) );
NOR2_X1 U21388 ( .A1(n19856), .A2(n2901), .ZN(n3000) );
NAND2_X1 U21389 ( .A1(n2994), .A2(n2995), .ZN(n14824) );
NOR2_X1 U21390 ( .A1(n2996), .A2(n2997), .ZN(n2994) );
NAND2_X1 U21391 ( .A1(n16445), .A2(n15994), .ZN(n2995) );
NOR2_X1 U21392 ( .A1(n19853), .A2(n16443), .ZN(n2996) );
INV_X1 U21393 ( .A(n21487), .ZN(n19936) );
INV_X1 U21394 ( .A(n22529), .ZN(n20900) );
INV_X1 U21395 ( .A(n22311), .ZN(n20896) );
NAND2_X1 U21396 ( .A1(n5134), .A2(n4051), .ZN(n15559) );
NAND2_X1 U21397 ( .A1(n5135), .A2(n15813), .ZN(n5134) );
NAND2_X1 U21398 ( .A1(n5136), .A2(n5137), .ZN(n5135) );
NOR2_X1 U21399 ( .A1(n20983), .A2(n5130), .ZN(n5136) );
NAND2_X1 U21400 ( .A1(n1927), .A2(n1928), .ZN(n15214) );
NAND2_X1 U21401 ( .A1(n16454), .A2(crash_dump_o_123_), .ZN(n1927) );
NAND2_X1 U21402 ( .A1(n16452), .A2(crash_dump_o_91_), .ZN(n1928) );
NAND2_X1 U21403 ( .A1(n1935), .A2(n1936), .ZN(n15184) );
NAND2_X1 U21404 ( .A1(n16456), .A2(crash_dump_o_121_), .ZN(n1935) );
NAND2_X1 U21405 ( .A1(n16452), .A2(crash_dump_o_89_), .ZN(n1936) );
NAND2_X1 U21406 ( .A1(n1939), .A2(n1940), .ZN(n15169) );
NAND2_X1 U21407 ( .A1(n16456), .A2(crash_dump_o_120_), .ZN(n1939) );
NAND2_X1 U21408 ( .A1(n16452), .A2(crash_dump_o_88_), .ZN(n1940) );
NAND2_X1 U21409 ( .A1(n1943), .A2(n1944), .ZN(n15154) );
NAND2_X1 U21410 ( .A1(n16457), .A2(crash_dump_o_119_), .ZN(n1943) );
NAND2_X1 U21411 ( .A1(n16452), .A2(crash_dump_o_87_), .ZN(n1944) );
NAND2_X1 U21412 ( .A1(n1947), .A2(n1948), .ZN(n15139) );
NAND2_X1 U21413 ( .A1(n16455), .A2(crash_dump_o_118_), .ZN(n1947) );
NAND2_X1 U21414 ( .A1(n16452), .A2(crash_dump_o_86_), .ZN(n1948) );
NAND2_X1 U21415 ( .A1(n1954), .A2(n1955), .ZN(n15124) );
NAND2_X1 U21416 ( .A1(n16457), .A2(crash_dump_o_116_), .ZN(n1954) );
NAND2_X1 U21417 ( .A1(n16452), .A2(crash_dump_o_84_), .ZN(n1955) );
NAND2_X1 U21418 ( .A1(n1961), .A2(n1962), .ZN(n15109) );
NAND2_X1 U21419 ( .A1(n16454), .A2(crash_dump_o_115_), .ZN(n1961) );
NAND2_X1 U21420 ( .A1(n16452), .A2(crash_dump_o_83_), .ZN(n1962) );
NAND2_X1 U21421 ( .A1(n1965), .A2(n1966), .ZN(n15092) );
NAND2_X1 U21422 ( .A1(n16455), .A2(crash_dump_o_114_), .ZN(n1965) );
NAND2_X1 U21423 ( .A1(n16452), .A2(crash_dump_o_82_), .ZN(n1966) );
NAND2_X1 U21424 ( .A1(n1973), .A2(n1974), .ZN(n15077) );
NAND2_X1 U21425 ( .A1(n16454), .A2(crash_dump_o_112_), .ZN(n1973) );
NAND2_X1 U21426 ( .A1(n16452), .A2(crash_dump_o_80_), .ZN(n1974) );
NAND2_X1 U21427 ( .A1(n1977), .A2(n1978), .ZN(n15062) );
NAND2_X1 U21428 ( .A1(n16456), .A2(crash_dump_o_111_), .ZN(n1977) );
NAND2_X1 U21429 ( .A1(n16452), .A2(crash_dump_o_79_), .ZN(n1978) );
NAND2_X1 U21430 ( .A1(n1981), .A2(n1982), .ZN(n15048) );
NAND2_X1 U21431 ( .A1(n16454), .A2(crash_dump_o_110_), .ZN(n1981) );
NAND2_X1 U21432 ( .A1(n16452), .A2(crash_dump_o_78_), .ZN(n1982) );
NAND2_X1 U21433 ( .A1(n1985), .A2(n1986), .ZN(n15033) );
NAND2_X1 U21434 ( .A1(n16456), .A2(crash_dump_o_109_), .ZN(n1985) );
NAND2_X1 U21435 ( .A1(n16452), .A2(crash_dump_o_77_), .ZN(n1986) );
NAND2_X1 U21436 ( .A1(n1989), .A2(n1990), .ZN(n15012) );
NAND2_X1 U21437 ( .A1(n16455), .A2(crash_dump_o_108_), .ZN(n1989) );
NAND2_X1 U21438 ( .A1(n16451), .A2(crash_dump_o_76_), .ZN(n1990) );
NAND2_X1 U21439 ( .A1(n1996), .A2(n1997), .ZN(n15003) );
NAND2_X1 U21440 ( .A1(n16457), .A2(crash_dump_o_106_), .ZN(n1996) );
NAND2_X1 U21441 ( .A1(n16451), .A2(crash_dump_o_74_), .ZN(n1997) );
NAND2_X1 U21442 ( .A1(n1969), .A2(n1970), .ZN(n14891) );
NAND2_X1 U21443 ( .A1(n16454), .A2(crash_dump_o_113_), .ZN(n1969) );
NAND2_X1 U21444 ( .A1(n16452), .A2(crash_dump_o_81_), .ZN(n1970) );
NAND2_X1 U21445 ( .A1(n3413), .A2(n3414), .ZN(n15781) );
NOR2_X1 U21446 ( .A1(n3415), .A2(n3416), .ZN(n3413) );
NAND2_X1 U21447 ( .A1(n16345), .A2(crash_dump_o_69_), .ZN(n3414) );
AND2_X1 U21448 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_5), .A2(n3396), .ZN(n3416) );
NAND2_X1 U21449 ( .A1(n3392), .A2(n3393), .ZN(n14990) );
NOR2_X1 U21450 ( .A1(n3394), .A2(n3395), .ZN(n3392) );
NAND2_X1 U21451 ( .A1(n16345), .A2(crash_dump_o_73_), .ZN(n3393) );
AND2_X1 U21452 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_9), .A2(n3396), .ZN(n3395) );
NAND2_X1 U21453 ( .A1(n3398), .A2(n3399), .ZN(n14976) );
NOR2_X1 U21454 ( .A1(n3400), .A2(n3401), .ZN(n3398) );
NAND2_X1 U21455 ( .A1(n16345), .A2(crash_dump_o_72_), .ZN(n3399) );
AND2_X1 U21456 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_8), .A2(n3396), .ZN(n3401) );
NAND2_X1 U21457 ( .A1(n3408), .A2(n3409), .ZN(n14962) );
NOR2_X1 U21458 ( .A1(n3410), .A2(n3411), .ZN(n3408) );
NAND2_X1 U21459 ( .A1(n16345), .A2(crash_dump_o_70_), .ZN(n3409) );
AND2_X1 U21460 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_6), .A2(n3396), .ZN(n3411) );
NAND2_X1 U21461 ( .A1(n3418), .A2(n3419), .ZN(n14949) );
NOR2_X1 U21462 ( .A1(n3420), .A2(n3421), .ZN(n3418) );
NAND2_X1 U21463 ( .A1(n16345), .A2(crash_dump_o_68_), .ZN(n3419) );
AND2_X1 U21464 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_4), .A2(n16432), .ZN(n3421) );
NAND2_X1 U21465 ( .A1(n3403), .A2(n3404), .ZN(n14925) );
NOR2_X1 U21466 ( .A1(n3405), .A2(n3406), .ZN(n3403) );
NAND2_X1 U21467 ( .A1(n16345), .A2(crash_dump_o_71_), .ZN(n3404) );
AND2_X1 U21468 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_7), .A2(n3396), .ZN(n3406) );
NAND2_X1 U21469 ( .A1(n1931), .A2(n1932), .ZN(n15199) );
NAND2_X1 U21470 ( .A1(n16455), .A2(crash_dump_o_122_), .ZN(n1931) );
NAND2_X1 U21471 ( .A1(n16453), .A2(crash_dump_o_90_), .ZN(n1932) );
NAND2_X1 U21472 ( .A1(n1889), .A2(n1890), .ZN(n14975) );
NAND2_X1 U21473 ( .A1(n16457), .A2(crash_dump_o_104_), .ZN(n1889) );
NAND2_X1 U21474 ( .A1(n16453), .A2(crash_dump_o_72_), .ZN(n1890) );
NAND2_X1 U21475 ( .A1(n1897), .A2(n1898), .ZN(n14961) );
NAND2_X1 U21476 ( .A1(n16457), .A2(crash_dump_o_102_), .ZN(n1897) );
NAND2_X1 U21477 ( .A1(n16453), .A2(crash_dump_o_70_), .ZN(n1898) );
NAND2_X1 U21478 ( .A1(n1893), .A2(n1894), .ZN(n14924) );
NAND2_X1 U21479 ( .A1(n16454), .A2(crash_dump_o_103_), .ZN(n1893) );
NAND2_X1 U21480 ( .A1(n16453), .A2(crash_dump_o_71_), .ZN(n1894) );
NAND2_X1 U21481 ( .A1(n1923), .A2(n1924), .ZN(n14875) );
NAND2_X1 U21482 ( .A1(n16455), .A2(crash_dump_o_124_), .ZN(n1923) );
NAND2_X1 U21483 ( .A1(n16453), .A2(crash_dump_o_92_), .ZN(n1924) );
NAND2_X1 U21484 ( .A1(n1919), .A2(n1920), .ZN(n14865) );
NAND2_X1 U21485 ( .A1(n16454), .A2(crash_dump_o_125_), .ZN(n1919) );
NAND2_X1 U21486 ( .A1(n16453), .A2(crash_dump_o_93_), .ZN(n1920) );
NAND2_X1 U21487 ( .A1(n2729), .A2(n2730), .ZN(n15623) );
NAND2_X1 U21488 ( .A1(n16454), .A2(n15894), .ZN(n2729) );
NAND2_X1 U21489 ( .A1(n16451), .A2(n2399), .ZN(n2730) );
NAND2_X1 U21490 ( .A1(n1883), .A2(n1884), .ZN(n14989) );
NAND2_X1 U21491 ( .A1(n16455), .A2(crash_dump_o_105_), .ZN(n1883) );
NAND2_X1 U21492 ( .A1(n16452), .A2(crash_dump_o_73_), .ZN(n1884) );
NAND2_X1 U21493 ( .A1(n3493), .A2(n3494), .ZN(n15762) );
NAND2_X1 U21494 ( .A1(n19883), .A2(crash_dump_o_65_), .ZN(n3494) );
NOR2_X1 U21495 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_add_243_A_1_), .A2(n3495), .ZN(n3493) );
AND2_X1 U21496 ( .A1(n3496), .A2(n16442), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_add_243_A_1_) );
NAND2_X1 U21497 ( .A1(n3544), .A2(n3545), .ZN(n15569) );
NAND2_X1 U21498 ( .A1(n16345), .A2(crash_dump_o_75_), .ZN(n3545) );
NOR2_X1 U21499 ( .A1(n3546), .A2(n3547), .ZN(n3544) );
AND2_X1 U21500 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_11), .A2(n3396), .ZN(n3546) );
NAND2_X1 U21501 ( .A1(n3488), .A2(n3489), .ZN(n15125) );
NAND2_X1 U21502 ( .A1(n19883), .A2(crash_dump_o_84_), .ZN(n3489) );
NOR2_X1 U21503 ( .A1(n3490), .A2(n3491), .ZN(n3488) );
AND2_X1 U21504 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_20), .A2(n16432), .ZN(n3490) );
NAND2_X1 U21505 ( .A1(n3504), .A2(n3505), .ZN(n15110) );
NAND2_X1 U21506 ( .A1(n16345), .A2(crash_dump_o_83_), .ZN(n3505) );
NOR2_X1 U21507 ( .A1(n3506), .A2(n3507), .ZN(n3504) );
AND2_X1 U21508 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_19), .A2(n16432), .ZN(n3507) );
NAND2_X1 U21509 ( .A1(n3509), .A2(n3510), .ZN(n15093) );
NAND2_X1 U21510 ( .A1(n19883), .A2(crash_dump_o_82_), .ZN(n3510) );
NOR2_X1 U21511 ( .A1(n3511), .A2(n3512), .ZN(n3509) );
AND2_X1 U21512 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_18), .A2(n16432), .ZN(n3512) );
NAND2_X1 U21513 ( .A1(n3519), .A2(n3520), .ZN(n15078) );
NAND2_X1 U21514 ( .A1(n16345), .A2(crash_dump_o_80_), .ZN(n3520) );
NOR2_X1 U21515 ( .A1(n3521), .A2(n3522), .ZN(n3519) );
AND2_X1 U21516 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_16), .A2(n3396), .ZN(n3521) );
NAND2_X1 U21517 ( .A1(n3524), .A2(n3525), .ZN(n15063) );
NAND2_X1 U21518 ( .A1(n19883), .A2(crash_dump_o_79_), .ZN(n3525) );
NOR2_X1 U21519 ( .A1(n3526), .A2(n3527), .ZN(n3524) );
AND2_X1 U21520 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_15), .A2(n3396), .ZN(n3527) );
NAND2_X1 U21521 ( .A1(n3529), .A2(n3530), .ZN(n15049) );
NAND2_X1 U21522 ( .A1(n16345), .A2(crash_dump_o_78_), .ZN(n3530) );
NOR2_X1 U21523 ( .A1(n3531), .A2(n3532), .ZN(n3529) );
AND2_X1 U21524 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_14), .A2(n3396), .ZN(n3532) );
NAND2_X1 U21525 ( .A1(n3534), .A2(n3535), .ZN(n15034) );
NAND2_X1 U21526 ( .A1(n19883), .A2(crash_dump_o_77_), .ZN(n3535) );
NOR2_X1 U21527 ( .A1(n3536), .A2(n3537), .ZN(n3534) );
AND2_X1 U21528 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_13), .A2(n3396), .ZN(n3537) );
NAND2_X1 U21529 ( .A1(n3539), .A2(n3540), .ZN(n15013) );
NAND2_X1 U21530 ( .A1(n16345), .A2(crash_dump_o_76_), .ZN(n3540) );
NOR2_X1 U21531 ( .A1(n3541), .A2(n3542), .ZN(n3539) );
AND2_X1 U21532 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_12), .A2(n3396), .ZN(n3542) );
NAND2_X1 U21533 ( .A1(n3549), .A2(n3550), .ZN(n15004) );
NAND2_X1 U21534 ( .A1(n19883), .A2(crash_dump_o_74_), .ZN(n3550) );
NOR2_X1 U21535 ( .A1(n3551), .A2(n3552), .ZN(n3549) );
AND2_X1 U21536 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_10), .A2(n3396), .ZN(n3552) );
NAND2_X1 U21537 ( .A1(n3514), .A2(n3515), .ZN(n14892) );
NAND2_X1 U21538 ( .A1(n16345), .A2(crash_dump_o_81_), .ZN(n3515) );
NOR2_X1 U21539 ( .A1(n3516), .A2(n3517), .ZN(n3514) );
AND2_X1 U21540 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_17), .A2(n16432), .ZN(n3517) );
NAND2_X1 U21541 ( .A1(n3428), .A2(n3429), .ZN(n15780) );
NAND2_X1 U21542 ( .A1(n19883), .A2(crash_dump_o_95_), .ZN(n3429) );
NOR2_X1 U21543 ( .A1(n3430), .A2(n3431), .ZN(n3428) );
AND2_X1 U21544 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_31), .A2(n16432), .ZN(n3431) );
NAND2_X1 U21545 ( .A1(n3433), .A2(n3434), .ZN(n15775) );
NAND2_X1 U21546 ( .A1(n19883), .A2(crash_dump_o_94_), .ZN(n3434) );
NOR2_X1 U21547 ( .A1(n3435), .A2(n3436), .ZN(n3433) );
AND2_X1 U21548 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_30), .A2(n3396), .ZN(n3436) );
NAND2_X1 U21549 ( .A1(n3483), .A2(n3484), .ZN(n15770) );
NAND2_X1 U21550 ( .A1(n19883), .A2(crash_dump_o_85_), .ZN(n3484) );
NOR2_X1 U21551 ( .A1(n3485), .A2(n3486), .ZN(n3483) );
AND2_X1 U21552 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_21), .A2(n16432), .ZN(n3486) );
NAND2_X1 U21553 ( .A1(n3453), .A2(n3454), .ZN(n15215) );
NAND2_X1 U21554 ( .A1(n19883), .A2(crash_dump_o_91_), .ZN(n3454) );
NOR2_X1 U21555 ( .A1(n3455), .A2(n3456), .ZN(n3453) );
AND2_X1 U21556 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_27), .A2(n16432), .ZN(n3455) );
NAND2_X1 U21557 ( .A1(n3458), .A2(n3459), .ZN(n15200) );
NAND2_X1 U21558 ( .A1(n19883), .A2(crash_dump_o_90_), .ZN(n3459) );
NOR2_X1 U21559 ( .A1(n3460), .A2(n3461), .ZN(n3458) );
AND2_X1 U21560 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_26), .A2(n16432), .ZN(n3461) );
NAND2_X1 U21561 ( .A1(n3463), .A2(n3464), .ZN(n15185) );
NAND2_X1 U21562 ( .A1(n19883), .A2(crash_dump_o_89_), .ZN(n3464) );
NOR2_X1 U21563 ( .A1(n3465), .A2(n3466), .ZN(n3463) );
AND2_X1 U21564 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_25), .A2(n16432), .ZN(n3465) );
NAND2_X1 U21565 ( .A1(n3468), .A2(n3469), .ZN(n15170) );
NAND2_X1 U21566 ( .A1(n16345), .A2(crash_dump_o_88_), .ZN(n3469) );
NOR2_X1 U21567 ( .A1(n3470), .A2(n3471), .ZN(n3468) );
AND2_X1 U21568 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_24), .A2(n16432), .ZN(n3471) );
NAND2_X1 U21569 ( .A1(n3473), .A2(n3474), .ZN(n15155) );
NAND2_X1 U21570 ( .A1(n19883), .A2(crash_dump_o_87_), .ZN(n3474) );
NOR2_X1 U21571 ( .A1(n3475), .A2(n3476), .ZN(n3473) );
AND2_X1 U21572 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_23), .A2(n16432), .ZN(n3476) );
NAND2_X1 U21573 ( .A1(n3478), .A2(n3479), .ZN(n15140) );
NAND2_X1 U21574 ( .A1(n16345), .A2(crash_dump_o_86_), .ZN(n3479) );
NOR2_X1 U21575 ( .A1(n3480), .A2(n3481), .ZN(n3478) );
AND2_X1 U21576 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_22), .A2(n16432), .ZN(n3481) );
NAND2_X1 U21577 ( .A1(n3423), .A2(n3424), .ZN(n14915) );
NAND2_X1 U21578 ( .A1(n19883), .A2(crash_dump_o_67_), .ZN(n3424) );
NOR2_X1 U21579 ( .A1(n3425), .A2(n3426), .ZN(n3423) );
AND2_X1 U21580 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_3), .A2(n16432), .ZN(n3426) );
NAND2_X1 U21581 ( .A1(n3438), .A2(n3439), .ZN(n14907) );
NAND2_X1 U21582 ( .A1(n16345), .A2(crash_dump_o_66_), .ZN(n3439) );
NOR2_X1 U21583 ( .A1(n3440), .A2(n3441), .ZN(n3438) );
AND2_X1 U21584 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_2), .A2(n3396), .ZN(n3441) );
NAND2_X1 U21585 ( .A1(n3448), .A2(n3449), .ZN(n14876) );
NAND2_X1 U21586 ( .A1(n19883), .A2(crash_dump_o_92_), .ZN(n3449) );
NOR2_X1 U21587 ( .A1(n3450), .A2(n3451), .ZN(n3448) );
AND2_X1 U21588 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_28), .A2(n16432), .ZN(n3450) );
NAND2_X1 U21589 ( .A1(n3443), .A2(n3444), .ZN(n14866) );
NAND2_X1 U21590 ( .A1(n16345), .A2(crash_dump_o_93_), .ZN(n3444) );
NOR2_X1 U21591 ( .A1(n3445), .A2(n3446), .ZN(n3443) );
AND2_X1 U21592 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_29), .A2(n3396), .ZN(n3446) );
NAND2_X1 U21593 ( .A1(n5543), .A2(n5544), .ZN(n15544) );
NAND2_X1 U21594 ( .A1(n5374), .A2(n15877), .ZN(n5544) );
NOR2_X1 U21595 ( .A1(n20999), .A2(n5545), .ZN(n5543) );
NOR2_X1 U21596 ( .A1(n5546), .A2(n5374), .ZN(n5545) );
NAND2_X1 U21597 ( .A1(n5533), .A2(n5534), .ZN(n15511) );
NAND2_X1 U21598 ( .A1(n5374), .A2(n15887), .ZN(n5534) );
NOR2_X1 U21599 ( .A1(n21001), .A2(n5535), .ZN(n5533) );
NOR2_X1 U21600 ( .A1(n5536), .A2(n5374), .ZN(n5535) );
NAND2_X1 U21601 ( .A1(n5419), .A2(n5420), .ZN(n15535) );
NAND2_X1 U21602 ( .A1(n5382), .A2(n16085), .ZN(n5420) );
NOR2_X1 U21603 ( .A1(n5421), .A2(n5422), .ZN(n5419) );
NOR2_X1 U21604 ( .A1(n20176), .A2(n16414), .ZN(n5422) );
NAND2_X1 U21605 ( .A1(n5438), .A2(n5439), .ZN(n15531) );
NAND2_X1 U21606 ( .A1(n5382), .A2(n16086), .ZN(n5439) );
NOR2_X1 U21607 ( .A1(n5440), .A2(n5441), .ZN(n5438) );
NOR2_X1 U21608 ( .A1(n20291), .A2(n5385), .ZN(n5441) );
NAND2_X1 U21609 ( .A1(n5442), .A2(n5443), .ZN(n15530) );
NAND2_X1 U21610 ( .A1(n16415), .A2(n16087), .ZN(n5443) );
NOR2_X1 U21611 ( .A1(n5444), .A2(n5445), .ZN(n5442) );
NOR2_X1 U21612 ( .A1(n20330), .A2(n16414), .ZN(n5445) );
NAND2_X1 U21613 ( .A1(n5451), .A2(n5452), .ZN(n15528) );
NAND2_X1 U21614 ( .A1(n5382), .A2(n16088), .ZN(n5452) );
NOR2_X1 U21615 ( .A1(n5453), .A2(n5454), .ZN(n5451) );
NOR2_X1 U21616 ( .A1(n20408), .A2(n5385), .ZN(n5454) );
NAND2_X1 U21617 ( .A1(n5455), .A2(n5456), .ZN(n15527) );
NAND2_X1 U21618 ( .A1(n16415), .A2(n16089), .ZN(n5456) );
NOR2_X1 U21619 ( .A1(n5457), .A2(n5458), .ZN(n5455) );
NOR2_X1 U21620 ( .A1(n20448), .A2(n16414), .ZN(n5458) );
NAND2_X1 U21621 ( .A1(n5459), .A2(n5460), .ZN(n15526) );
NAND2_X1 U21622 ( .A1(n5382), .A2(n16090), .ZN(n5460) );
NOR2_X1 U21623 ( .A1(n5461), .A2(n5462), .ZN(n5459) );
NOR2_X1 U21624 ( .A1(n20488), .A2(n5385), .ZN(n5462) );
NAND2_X1 U21625 ( .A1(n5463), .A2(n5464), .ZN(n15525) );
NAND2_X1 U21626 ( .A1(n16415), .A2(n16091), .ZN(n5464) );
NOR2_X1 U21627 ( .A1(n5465), .A2(n5466), .ZN(n5463) );
NOR2_X1 U21628 ( .A1(n20528), .A2(n16414), .ZN(n5466) );
NAND2_X1 U21629 ( .A1(n5467), .A2(n5468), .ZN(n15524) );
NAND2_X1 U21630 ( .A1(n5382), .A2(n16092), .ZN(n5468) );
NOR2_X1 U21631 ( .A1(n5469), .A2(n5470), .ZN(n5467) );
NOR2_X1 U21632 ( .A1(n20568), .A2(n5385), .ZN(n5470) );
NAND2_X1 U21633 ( .A1(n5471), .A2(n5472), .ZN(n15523) );
NAND2_X1 U21634 ( .A1(n5382), .A2(n16120), .ZN(n5472) );
NOR2_X1 U21635 ( .A1(n5473), .A2(n5474), .ZN(n5471) );
NOR2_X1 U21636 ( .A1(n20756), .A2(n16414), .ZN(n5474) );
NAND2_X1 U21637 ( .A1(n5505), .A2(n5506), .ZN(n15516) );
NAND2_X1 U21638 ( .A1(n5382), .A2(n16093), .ZN(n5506) );
NOR2_X1 U21639 ( .A1(n5507), .A2(n5508), .ZN(n5505) );
NOR2_X1 U21640 ( .A1(n20699), .A2(n5385), .ZN(n5508) );
NAND2_X1 U21641 ( .A1(n5509), .A2(n5510), .ZN(n15515) );
NAND2_X1 U21642 ( .A1(n5382), .A2(n16094), .ZN(n5510) );
NOR2_X1 U21643 ( .A1(n5511), .A2(n5512), .ZN(n5509) );
NOR2_X1 U21644 ( .A1(n20703), .A2(n16414), .ZN(n5512) );
NAND2_X1 U21645 ( .A1(n4110), .A2(n4111), .ZN(n15497) );
NAND2_X1 U21646 ( .A1(n4061), .A2(n16095), .ZN(n4111) );
NOR2_X1 U21647 ( .A1(n4113), .A2(n4114), .ZN(n4110) );
NOR2_X1 U21648 ( .A1(n20767), .A2(n4066), .ZN(n4114) );
NAND2_X1 U21649 ( .A1(n4122), .A2(n4123), .ZN(n15495) );
NAND2_X1 U21650 ( .A1(n4061), .A2(n16096), .ZN(n4123) );
NOR2_X1 U21651 ( .A1(n4125), .A2(n4126), .ZN(n4122) );
NOR2_X1 U21652 ( .A1(n20770), .A2(n16426), .ZN(n4126) );
NAND2_X1 U21653 ( .A1(n4128), .A2(n4129), .ZN(n15494) );
NAND2_X1 U21654 ( .A1(n4061), .A2(n16097), .ZN(n4129) );
NOR2_X1 U21655 ( .A1(n4131), .A2(n4132), .ZN(n4128) );
NOR2_X1 U21656 ( .A1(n20773), .A2(n4066), .ZN(n4132) );
NAND2_X1 U21657 ( .A1(n4134), .A2(n4135), .ZN(n15493) );
NAND2_X1 U21658 ( .A1(n4061), .A2(n16098), .ZN(n4135) );
NOR2_X1 U21659 ( .A1(n4137), .A2(n4138), .ZN(n4134) );
NOR2_X1 U21660 ( .A1(n20776), .A2(n16426), .ZN(n4138) );
NAND2_X1 U21661 ( .A1(n4140), .A2(n4141), .ZN(n15492) );
NAND2_X1 U21662 ( .A1(n4061), .A2(n16099), .ZN(n4141) );
NOR2_X1 U21663 ( .A1(n4143), .A2(n4144), .ZN(n4140) );
NOR2_X1 U21664 ( .A1(n20779), .A2(n4066), .ZN(n4144) );
NAND2_X1 U21665 ( .A1(n4146), .A2(n4147), .ZN(n15491) );
NAND2_X1 U21666 ( .A1(n4061), .A2(n16100), .ZN(n4147) );
NOR2_X1 U21667 ( .A1(n4149), .A2(n4150), .ZN(n4146) );
NOR2_X1 U21668 ( .A1(n20782), .A2(n16426), .ZN(n4150) );
NAND2_X1 U21669 ( .A1(n4152), .A2(n4153), .ZN(n15490) );
NAND2_X1 U21670 ( .A1(n4061), .A2(n16101), .ZN(n4153) );
NOR2_X1 U21671 ( .A1(n4155), .A2(n4156), .ZN(n4152) );
NOR2_X1 U21672 ( .A1(n20785), .A2(n4066), .ZN(n4156) );
NAND2_X1 U21673 ( .A1(n4158), .A2(n4159), .ZN(n15489) );
NAND2_X1 U21674 ( .A1(n4061), .A2(n16102), .ZN(n4159) );
NOR2_X1 U21675 ( .A1(n4161), .A2(n4162), .ZN(n4158) );
NOR2_X1 U21676 ( .A1(n20788), .A2(n16426), .ZN(n4162) );
NAND2_X1 U21677 ( .A1(n4164), .A2(n4165), .ZN(n15488) );
NAND2_X1 U21678 ( .A1(n4061), .A2(n16103), .ZN(n4165) );
NOR2_X1 U21679 ( .A1(n4167), .A2(n4168), .ZN(n4164) );
NOR2_X1 U21680 ( .A1(n20791), .A2(n4066), .ZN(n4168) );
NAND2_X1 U21681 ( .A1(n4170), .A2(n4171), .ZN(n15487) );
NAND2_X1 U21682 ( .A1(n16427), .A2(n16104), .ZN(n4171) );
NOR2_X1 U21683 ( .A1(n4173), .A2(n4174), .ZN(n4170) );
NOR2_X1 U21684 ( .A1(n20794), .A2(n16426), .ZN(n4174) );
NAND2_X1 U21685 ( .A1(n4176), .A2(n4177), .ZN(n15486) );
NAND2_X1 U21686 ( .A1(n4061), .A2(n16105), .ZN(n4177) );
NOR2_X1 U21687 ( .A1(n4179), .A2(n4180), .ZN(n4176) );
NOR2_X1 U21688 ( .A1(n20797), .A2(n4066), .ZN(n4180) );
NAND2_X1 U21689 ( .A1(n4188), .A2(n4189), .ZN(n15484) );
NAND2_X1 U21690 ( .A1(n16427), .A2(n16106), .ZN(n4189) );
NOR2_X1 U21691 ( .A1(n4191), .A2(n4192), .ZN(n4188) );
NOR2_X1 U21692 ( .A1(n20800), .A2(n4066), .ZN(n4192) );
NAND2_X1 U21693 ( .A1(n4194), .A2(n4195), .ZN(n15483) );
NAND2_X1 U21694 ( .A1(n16427), .A2(n16107), .ZN(n4195) );
NOR2_X1 U21695 ( .A1(n4197), .A2(n4198), .ZN(n4194) );
NOR2_X1 U21696 ( .A1(n20803), .A2(n4066), .ZN(n4198) );
NAND2_X1 U21697 ( .A1(n4200), .A2(n4201), .ZN(n15482) );
NAND2_X1 U21698 ( .A1(n16427), .A2(n16108), .ZN(n4201) );
NOR2_X1 U21699 ( .A1(n4203), .A2(n4204), .ZN(n4200) );
NOR2_X1 U21700 ( .A1(n20806), .A2(n4066), .ZN(n4204) );
NAND2_X1 U21701 ( .A1(n4206), .A2(n4207), .ZN(n15481) );
NAND2_X1 U21702 ( .A1(n16427), .A2(n16109), .ZN(n4207) );
NOR2_X1 U21703 ( .A1(n4209), .A2(n4210), .ZN(n4206) );
NOR2_X1 U21704 ( .A1(n20809), .A2(n16426), .ZN(n4210) );
NAND2_X1 U21705 ( .A1(n4212), .A2(n4213), .ZN(n15480) );
NAND2_X1 U21706 ( .A1(n16427), .A2(n16110), .ZN(n4213) );
NOR2_X1 U21707 ( .A1(n4215), .A2(n4216), .ZN(n4212) );
NOR2_X1 U21708 ( .A1(n20811), .A2(n4066), .ZN(n4216) );
NAND2_X1 U21709 ( .A1(n4218), .A2(n4219), .ZN(n15479) );
NAND2_X1 U21710 ( .A1(n16427), .A2(n16111), .ZN(n4219) );
NOR2_X1 U21711 ( .A1(n4221), .A2(n4222), .ZN(n4218) );
NOR2_X1 U21712 ( .A1(n20813), .A2(n16426), .ZN(n4222) );
NAND2_X1 U21713 ( .A1(n4224), .A2(n4225), .ZN(n15478) );
NAND2_X1 U21714 ( .A1(n16427), .A2(n16112), .ZN(n4225) );
NOR2_X1 U21715 ( .A1(n4227), .A2(n4228), .ZN(n4224) );
NOR2_X1 U21716 ( .A1(n20815), .A2(n4066), .ZN(n4228) );
NAND2_X1 U21717 ( .A1(n4230), .A2(n4231), .ZN(n15477) );
NAND2_X1 U21718 ( .A1(n16427), .A2(n16113), .ZN(n4231) );
NOR2_X1 U21719 ( .A1(n4233), .A2(n4234), .ZN(n4230) );
NOR2_X1 U21720 ( .A1(n20817), .A2(n16426), .ZN(n4234) );
NAND2_X1 U21721 ( .A1(n5370), .A2(n5371), .ZN(n15409) );
NAND2_X1 U21722 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_0), .ZN(n5371) );
NAND2_X1 U21723 ( .A1(n5278), .A2(n16114), .ZN(n5370) );
NAND2_X1 U21724 ( .A1(n2934), .A2(n2935), .ZN(n14850) );
NAND2_X1 U21725 ( .A1(n2897), .A2(n15934), .ZN(n2935) );
NOR2_X1 U21726 ( .A1(n2936), .A2(n2937), .ZN(n2934) );
NOR2_X1 U21727 ( .A1(n20748), .A2(n2901), .ZN(n2936) );
NAND2_X1 U21728 ( .A1(n2922), .A2(n2923), .ZN(n14848) );
NAND2_X1 U21729 ( .A1(n2897), .A2(n15935), .ZN(n2923) );
NOR2_X1 U21730 ( .A1(n2924), .A2(n2925), .ZN(n2922) );
NOR2_X1 U21731 ( .A1(n20742), .A2(n2901), .ZN(n2924) );
NAND2_X1 U21732 ( .A1(n2918), .A2(n2919), .ZN(n14846) );
NAND2_X1 U21733 ( .A1(n2897), .A2(n15936), .ZN(n2919) );
NOR2_X1 U21734 ( .A1(n2920), .A2(n2921), .ZN(n2918) );
NOR2_X1 U21735 ( .A1(n20737), .A2(n16443), .ZN(n2920) );
NAND2_X1 U21736 ( .A1(n2914), .A2(n2915), .ZN(n14844) );
NAND2_X1 U21737 ( .A1(n2897), .A2(n16007), .ZN(n2915) );
NOR2_X1 U21738 ( .A1(n2916), .A2(n2917), .ZN(n2914) );
NOR2_X1 U21739 ( .A1(n20731), .A2(n2901), .ZN(n2916) );
NAND2_X1 U21740 ( .A1(n2910), .A2(n2911), .ZN(n14842) );
NAND2_X1 U21741 ( .A1(n2897), .A2(n15997), .ZN(n2911) );
NOR2_X1 U21742 ( .A1(n2912), .A2(n2913), .ZN(n2910) );
NOR2_X1 U21743 ( .A1(n20726), .A2(n2901), .ZN(n2912) );
NAND2_X1 U21744 ( .A1(n2906), .A2(n2907), .ZN(n14840) );
NAND2_X1 U21745 ( .A1(n2897), .A2(n16002), .ZN(n2907) );
NOR2_X1 U21746 ( .A1(n2908), .A2(n2909), .ZN(n2906) );
NOR2_X1 U21747 ( .A1(n20720), .A2(n16443), .ZN(n2908) );
NAND2_X1 U21748 ( .A1(n2902), .A2(n2903), .ZN(n14838) );
NAND2_X1 U21749 ( .A1(n16445), .A2(n15998), .ZN(n2903) );
NOR2_X1 U21750 ( .A1(n2904), .A2(n2905), .ZN(n2902) );
NOR2_X1 U21751 ( .A1(n19871), .A2(n16443), .ZN(n2904) );
NAND2_X1 U21752 ( .A1(n2895), .A2(n2896), .ZN(n14836) );
NAND2_X1 U21753 ( .A1(n2897), .A2(n15999), .ZN(n2896) );
NOR2_X1 U21754 ( .A1(n2898), .A2(n2899), .ZN(n2895) );
NOR2_X1 U21755 ( .A1(n19868), .A2(n2901), .ZN(n2898) );
NAND2_X1 U21756 ( .A1(n2986), .A2(n2987), .ZN(n14820) );
NAND2_X1 U21757 ( .A1(n2897), .A2(n15995), .ZN(n2987) );
NOR2_X1 U21758 ( .A1(n2988), .A2(n2989), .ZN(n2986) );
NOR2_X1 U21759 ( .A1(n19848), .A2(n16443), .ZN(n2988) );
NAND2_X1 U21760 ( .A1(n2982), .A2(n2983), .ZN(n14818) );
NAND2_X1 U21761 ( .A1(n16445), .A2(n15986), .ZN(n2983) );
NOR2_X1 U21762 ( .A1(n2984), .A2(n2985), .ZN(n2982) );
NOR2_X1 U21763 ( .A1(n19846), .A2(n16443), .ZN(n2984) );
NAND2_X1 U21764 ( .A1(n2978), .A2(n2979), .ZN(n14816) );
NAND2_X1 U21765 ( .A1(n2897), .A2(n15987), .ZN(n2979) );
NOR2_X1 U21766 ( .A1(n2980), .A2(n2981), .ZN(n2978) );
NOR2_X1 U21767 ( .A1(n19843), .A2(n16443), .ZN(n2980) );
NAND2_X1 U21768 ( .A1(n2970), .A2(n2971), .ZN(n14812) );
NAND2_X1 U21769 ( .A1(n16445), .A2(n15988), .ZN(n2971) );
NOR2_X1 U21770 ( .A1(n2972), .A2(n2973), .ZN(n2970) );
NOR2_X1 U21771 ( .A1(n19838), .A2(n16443), .ZN(n2972) );
NAND2_X1 U21772 ( .A1(n2966), .A2(n2967), .ZN(n14810) );
NAND2_X1 U21773 ( .A1(n2897), .A2(n15989), .ZN(n2967) );
NOR2_X1 U21774 ( .A1(n2968), .A2(n2969), .ZN(n2966) );
NOR2_X1 U21775 ( .A1(n19836), .A2(n2901), .ZN(n2968) );
NAND2_X1 U21776 ( .A1(n2962), .A2(n2963), .ZN(n14808) );
NAND2_X1 U21777 ( .A1(n16445), .A2(n15990), .ZN(n2963) );
NOR2_X1 U21778 ( .A1(n2964), .A2(n2965), .ZN(n2962) );
NOR2_X1 U21779 ( .A1(n19833), .A2(n2901), .ZN(n2964) );
NAND2_X1 U21780 ( .A1(n2958), .A2(n2959), .ZN(n14806) );
NAND2_X1 U21781 ( .A1(n2897), .A2(n15983), .ZN(n2959) );
NOR2_X1 U21782 ( .A1(n2960), .A2(n2961), .ZN(n2958) );
NOR2_X1 U21783 ( .A1(n19831), .A2(n16443), .ZN(n2960) );
NAND2_X1 U21784 ( .A1(n2950), .A2(n2951), .ZN(n14802) );
NAND2_X1 U21785 ( .A1(n16445), .A2(n15984), .ZN(n2951) );
NOR2_X1 U21786 ( .A1(n2952), .A2(n2953), .ZN(n2950) );
NOR2_X1 U21787 ( .A1(n19826), .A2(n16443), .ZN(n2952) );
NAND2_X1 U21788 ( .A1(n2938), .A2(n2939), .ZN(n14796) );
NAND2_X1 U21789 ( .A1(n16445), .A2(n15985), .ZN(n2939) );
NOR2_X1 U21790 ( .A1(n2940), .A2(n2941), .ZN(n2938) );
NOR2_X1 U21791 ( .A1(n19818), .A2(n16443), .ZN(n2940) );
NAND2_X1 U21792 ( .A1(n2930), .A2(n2931), .ZN(n14794) );
NAND2_X1 U21793 ( .A1(n2897), .A2(n15980), .ZN(n2931) );
NOR2_X1 U21794 ( .A1(n2932), .A2(n2933), .ZN(n2930) );
NOR2_X1 U21795 ( .A1(n19815), .A2(n16443), .ZN(n2932) );
NAND2_X1 U21796 ( .A1(n2926), .A2(n2927), .ZN(n14792) );
NAND2_X1 U21797 ( .A1(n16445), .A2(n15981), .ZN(n2927) );
NOR2_X1 U21798 ( .A1(n2928), .A2(n2929), .ZN(n2926) );
NOR2_X1 U21799 ( .A1(n19813), .A2(n2901), .ZN(n2928) );
NAND2_X1 U21800 ( .A1(n1504), .A2(n1505), .ZN(n15313) );
NAND2_X1 U21801 ( .A1(n1507), .A2(n15923), .ZN(n1504) );
NAND2_X1 U21802 ( .A1(n19963), .A2(alu_adder_result_ex_1), .ZN(n1505) );
NAND2_X1 U21803 ( .A1(n1655), .A2(n1656), .ZN(n15281) );
NAND2_X1 U21804 ( .A1(n16461), .A2(crash_dump_o_33_), .ZN(n1655) );
NAND2_X1 U21805 ( .A1(n1657), .A2(alu_adder_result_ex_1), .ZN(n1656) );
NAND2_X1 U21806 ( .A1(n1586), .A2(n1587), .ZN(n15315) );
NAND2_X1 U21807 ( .A1(n1507), .A2(n16115), .ZN(n1586) );
NAND2_X1 U21808 ( .A1(n1564), .A2(n19963), .ZN(n1587) );
NAND2_X1 U21809 ( .A1(n1625), .A2(n1626), .ZN(n15311) );
NAND2_X1 U21810 ( .A1(n16461), .A2(crash_dump_o_63_), .ZN(n1626) );
NAND2_X1 U21811 ( .A1(data_addr_o_31_), .A2(n1606), .ZN(n1625) );
NAND2_X1 U21812 ( .A1(n1628), .A2(n1629), .ZN(n15310) );
NAND2_X1 U21813 ( .A1(n16461), .A2(crash_dump_o_62_), .ZN(n1629) );
NAND2_X1 U21814 ( .A1(data_addr_o_30_), .A2(n1606), .ZN(n1628) );
NAND2_X1 U21815 ( .A1(n1650), .A2(n1651), .ZN(n15301) );
NAND2_X1 U21816 ( .A1(n16461), .A2(crash_dump_o_53_), .ZN(n1651) );
NAND2_X1 U21817 ( .A1(data_addr_o_21_), .A2(n1606), .ZN(n1650) );
NAND2_X1 U21818 ( .A1(n1667), .A2(n1668), .ZN(n15295) );
NAND2_X1 U21819 ( .A1(n16461), .A2(crash_dump_o_47_), .ZN(n1668) );
NAND2_X1 U21820 ( .A1(data_addr_o_15_), .A2(n1606), .ZN(n1667) );
NAND2_X1 U21821 ( .A1(n1670), .A2(n1671), .ZN(n15294) );
NAND2_X1 U21822 ( .A1(n16461), .A2(crash_dump_o_46_), .ZN(n1671) );
NAND2_X1 U21823 ( .A1(data_addr_o_14_), .A2(n16460), .ZN(n1670) );
NAND2_X1 U21824 ( .A1(n1673), .A2(n1674), .ZN(n15293) );
NAND2_X1 U21825 ( .A1(n16461), .A2(crash_dump_o_45_), .ZN(n1674) );
NAND2_X1 U21826 ( .A1(data_addr_o_13_), .A2(n16460), .ZN(n1673) );
NAND2_X1 U21827 ( .A1(n1676), .A2(n1677), .ZN(n15292) );
NAND2_X1 U21828 ( .A1(n16461), .A2(crash_dump_o_44_), .ZN(n1677) );
NAND2_X1 U21829 ( .A1(data_addr_o_12_), .A2(n1606), .ZN(n1676) );
NAND2_X1 U21830 ( .A1(n1679), .A2(n1680), .ZN(n15291) );
NAND2_X1 U21831 ( .A1(n16461), .A2(crash_dump_o_43_), .ZN(n1680) );
NAND2_X1 U21832 ( .A1(data_addr_o_11_), .A2(n16460), .ZN(n1679) );
NAND2_X1 U21833 ( .A1(n1682), .A2(n1683), .ZN(n15290) );
NAND2_X1 U21834 ( .A1(n16461), .A2(crash_dump_o_42_), .ZN(n1683) );
NAND2_X1 U21835 ( .A1(data_addr_o_10_), .A2(n1606), .ZN(n1682) );
NAND2_X1 U21836 ( .A1(n1602), .A2(n1603), .ZN(n15289) );
NAND2_X1 U21837 ( .A1(n16461), .A2(crash_dump_o_41_), .ZN(n1603) );
NAND2_X1 U21838 ( .A1(data_addr_o_9_), .A2(n1606), .ZN(n1602) );
NAND2_X1 U21839 ( .A1(n1607), .A2(n1608), .ZN(n15288) );
NAND2_X1 U21840 ( .A1(n16461), .A2(crash_dump_o_40_), .ZN(n1608) );
NAND2_X1 U21841 ( .A1(data_addr_o_8_), .A2(n16460), .ZN(n1607) );
NAND2_X1 U21842 ( .A1(n1610), .A2(n1611), .ZN(n15287) );
NAND2_X1 U21843 ( .A1(n16461), .A2(crash_dump_o_39_), .ZN(n1611) );
NAND2_X1 U21844 ( .A1(data_addr_o_7_), .A2(n16460), .ZN(n1610) );
NAND2_X1 U21845 ( .A1(n1613), .A2(n1614), .ZN(n15286) );
NAND2_X1 U21846 ( .A1(n16461), .A2(crash_dump_o_38_), .ZN(n1614) );
NAND2_X1 U21847 ( .A1(data_addr_o_6_), .A2(n1606), .ZN(n1613) );
NAND2_X1 U21848 ( .A1(n1616), .A2(n1617), .ZN(n15285) );
NAND2_X1 U21849 ( .A1(n16461), .A2(crash_dump_o_37_), .ZN(n1617) );
NAND2_X1 U21850 ( .A1(data_addr_o_5_), .A2(n1606), .ZN(n1616) );
NAND2_X1 U21851 ( .A1(n1619), .A2(n1620), .ZN(n15284) );
NAND2_X1 U21852 ( .A1(n16461), .A2(crash_dump_o_36_), .ZN(n1620) );
NAND2_X1 U21853 ( .A1(data_addr_o_4_), .A2(n1606), .ZN(n1619) );
NAND2_X1 U21854 ( .A1(n1622), .A2(n1623), .ZN(n15283) );
NAND2_X1 U21855 ( .A1(n16461), .A2(crash_dump_o_35_), .ZN(n1623) );
NAND2_X1 U21856 ( .A1(data_addr_o_3_), .A2(n16460), .ZN(n1622) );
NAND2_X1 U21857 ( .A1(n1631), .A2(n1632), .ZN(n15282) );
NAND2_X1 U21858 ( .A1(n16461), .A2(crash_dump_o_34_), .ZN(n1632) );
NAND2_X1 U21859 ( .A1(data_addr_o_2_), .A2(n1606), .ZN(n1631) );
NAND2_X1 U21860 ( .A1(n3636), .A2(n3637), .ZN(n14851) );
NAND2_X1 U21861 ( .A1(n16431), .A2(n15937), .ZN(n3637) );
NAND2_X1 U21862 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_2), .A2(n3611), .ZN(n3636) );
NAND2_X1 U21863 ( .A1(n21375), .A2(n21374), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_2) );
NAND2_X1 U21864 ( .A1(n3627), .A2(n3628), .ZN(n14849) );
NAND2_X1 U21865 ( .A1(n16431), .A2(n16126), .ZN(n3628) );
NAND2_X1 U21866 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_3), .A2(n3611), .ZN(n3627) );
NAND2_X1 U21867 ( .A1(n21386), .A2(n21385), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_3) );
NAND2_X1 U21868 ( .A1(n3624), .A2(n3625), .ZN(n14847) );
NAND2_X1 U21869 ( .A1(n16431), .A2(n15938), .ZN(n3625) );
NAND2_X1 U21870 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_4), .A2(n3611), .ZN(n3624) );
NAND2_X1 U21871 ( .A1(n21388), .A2(n21387), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_4) );
NAND2_X1 U21872 ( .A1(n3621), .A2(n3622), .ZN(n14845) );
NAND2_X1 U21873 ( .A1(n16431), .A2(n15939), .ZN(n3622) );
NAND2_X1 U21874 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_5), .A2(n3611), .ZN(n3621) );
NAND2_X1 U21875 ( .A1(n21392), .A2(n21391), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_5) );
NAND2_X1 U21876 ( .A1(n3618), .A2(n3619), .ZN(n14843) );
NAND2_X1 U21877 ( .A1(n16430), .A2(n15940), .ZN(n3619) );
NAND2_X1 U21878 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_6), .A2(n3611), .ZN(n3618) );
NAND2_X1 U21879 ( .A1(n21394), .A2(n21393), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_6) );
NAND2_X1 U21880 ( .A1(n3615), .A2(n3616), .ZN(n14841) );
NAND2_X1 U21881 ( .A1(n16430), .A2(n15941), .ZN(n3616) );
NAND2_X1 U21882 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_7), .A2(n16429), .ZN(n3615) );
NAND2_X1 U21883 ( .A1(n21398), .A2(n21397), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_7) );
NAND2_X1 U21884 ( .A1(n3612), .A2(n3613), .ZN(n14839) );
NAND2_X1 U21885 ( .A1(n16431), .A2(n15942), .ZN(n3613) );
NAND2_X1 U21886 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_8), .A2(n16429), .ZN(n3612) );
NAND2_X1 U21887 ( .A1(n21400), .A2(n21399), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_8) );
NAND2_X1 U21888 ( .A1(n3607), .A2(n3608), .ZN(n14837) );
NAND2_X1 U21889 ( .A1(n16430), .A2(n15943), .ZN(n3608) );
NAND2_X1 U21890 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_9), .A2(n3611), .ZN(n3607) );
NAND2_X1 U21891 ( .A1(n21404), .A2(n21403), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_9) );
NAND2_X1 U21892 ( .A1(n3696), .A2(n3697), .ZN(n14835) );
NAND2_X1 U21893 ( .A1(n16431), .A2(n15944), .ZN(n3697) );
NAND2_X1 U21894 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_10), .A2(n3611), .ZN(n3696) );
NAND2_X1 U21895 ( .A1(n21307), .A2(n21306), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_10) );
NAND2_X1 U21896 ( .A1(n3693), .A2(n3694), .ZN(n14833) );
NAND2_X1 U21897 ( .A1(n16431), .A2(n15945), .ZN(n3694) );
NAND2_X1 U21898 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_11), .A2(n16429), .ZN(n3693) );
NAND2_X1 U21899 ( .A1(n21310), .A2(n21309), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_11) );
NAND2_X1 U21900 ( .A1(n3690), .A2(n3691), .ZN(n14831) );
NAND2_X1 U21901 ( .A1(n16431), .A2(n15946), .ZN(n3691) );
NAND2_X1 U21902 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_12), .A2(n16429), .ZN(n3690) );
NAND2_X1 U21903 ( .A1(n21314), .A2(n21313), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_12) );
NAND2_X1 U21904 ( .A1(n3687), .A2(n3688), .ZN(n14829) );
NAND2_X1 U21905 ( .A1(n16430), .A2(n15947), .ZN(n3688) );
NAND2_X1 U21906 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_13), .A2(n16429), .ZN(n3687) );
NAND2_X1 U21907 ( .A1(n21317), .A2(n21316), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_13) );
NAND2_X1 U21908 ( .A1(n3684), .A2(n3685), .ZN(n14827) );
NAND2_X1 U21909 ( .A1(n16431), .A2(n15948), .ZN(n3685) );
NAND2_X1 U21910 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_14), .A2(n16429), .ZN(n3684) );
NAND2_X1 U21911 ( .A1(n21321), .A2(n21320), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_14) );
NAND2_X1 U21912 ( .A1(n3681), .A2(n3682), .ZN(n14825) );
NAND2_X1 U21913 ( .A1(n16430), .A2(n15949), .ZN(n3682) );
NAND2_X1 U21914 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_15), .A2(n3611), .ZN(n3681) );
NAND2_X1 U21915 ( .A1(n21324), .A2(n21323), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_15) );
NAND2_X1 U21916 ( .A1(n3678), .A2(n3679), .ZN(n14823) );
NAND2_X1 U21917 ( .A1(n16430), .A2(n15950), .ZN(n3679) );
NAND2_X1 U21918 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_16), .A2(n3611), .ZN(n3678) );
NAND2_X1 U21919 ( .A1(n21328), .A2(n21327), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_16) );
NAND2_X1 U21920 ( .A1(n3675), .A2(n3676), .ZN(n14821) );
NAND2_X1 U21921 ( .A1(n16430), .A2(n15951), .ZN(n3676) );
NAND2_X1 U21922 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_17), .A2(n3611), .ZN(n3675) );
NAND2_X1 U21923 ( .A1(n21331), .A2(n21330), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_17) );
NAND2_X1 U21924 ( .A1(n3672), .A2(n3673), .ZN(n14819) );
NAND2_X1 U21925 ( .A1(n16430), .A2(n15952), .ZN(n3673) );
NAND2_X1 U21926 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_18), .A2(n3611), .ZN(n3672) );
NAND2_X1 U21927 ( .A1(n21335), .A2(n21334), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_18) );
NAND2_X1 U21928 ( .A1(n3669), .A2(n3670), .ZN(n14817) );
NAND2_X1 U21929 ( .A1(n16431), .A2(n15953), .ZN(n3670) );
NAND2_X1 U21930 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_19), .A2(n16429), .ZN(n3669) );
NAND2_X1 U21931 ( .A1(n21338), .A2(n21337), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_19) );
NAND2_X1 U21932 ( .A1(n3666), .A2(n3667), .ZN(n14815) );
NAND2_X1 U21933 ( .A1(n16430), .A2(n15954), .ZN(n3667) );
NAND2_X1 U21934 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_20), .A2(n16429), .ZN(n3666) );
NAND2_X1 U21935 ( .A1(n21342), .A2(n21341), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_20) );
NAND2_X1 U21936 ( .A1(n3663), .A2(n3664), .ZN(n14813) );
NAND2_X1 U21937 ( .A1(n16431), .A2(n15955), .ZN(n3664) );
NAND2_X1 U21938 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_21), .A2(n3611), .ZN(n3663) );
NAND2_X1 U21939 ( .A1(n21345), .A2(n21344), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_21) );
NAND2_X1 U21940 ( .A1(n3660), .A2(n3661), .ZN(n14811) );
NAND2_X1 U21941 ( .A1(n16430), .A2(n15956), .ZN(n3661) );
NAND2_X1 U21942 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_22), .A2(n16429), .ZN(n3660) );
NAND2_X1 U21943 ( .A1(n21349), .A2(n21348), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_22) );
NAND2_X1 U21944 ( .A1(n3657), .A2(n3658), .ZN(n14809) );
NAND2_X1 U21945 ( .A1(n16430), .A2(n15957), .ZN(n3658) );
NAND2_X1 U21946 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_23), .A2(n16429), .ZN(n3657) );
NAND2_X1 U21947 ( .A1(n21352), .A2(n21351), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_23) );
NAND2_X1 U21948 ( .A1(n3654), .A2(n3655), .ZN(n14807) );
NAND2_X1 U21949 ( .A1(n16430), .A2(n15958), .ZN(n3655) );
NAND2_X1 U21950 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_24), .A2(n16429), .ZN(n3654) );
NAND2_X1 U21951 ( .A1(n21356), .A2(n21355), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_24) );
NAND2_X1 U21952 ( .A1(n3651), .A2(n3652), .ZN(n14805) );
NAND2_X1 U21953 ( .A1(n16431), .A2(n15959), .ZN(n3652) );
NAND2_X1 U21954 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_25), .A2(n16429), .ZN(n3651) );
NAND2_X1 U21955 ( .A1(n21359), .A2(n21358), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_25) );
NAND2_X1 U21956 ( .A1(n3648), .A2(n3649), .ZN(n14803) );
NAND2_X1 U21957 ( .A1(n16430), .A2(n15960), .ZN(n3649) );
NAND2_X1 U21958 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_26), .A2(n3611), .ZN(n3648) );
NAND2_X1 U21959 ( .A1(n21363), .A2(n21362), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_26) );
NAND2_X1 U21960 ( .A1(n3645), .A2(n3646), .ZN(n14801) );
NAND2_X1 U21961 ( .A1(n16430), .A2(n15961), .ZN(n3646) );
NAND2_X1 U21962 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_27), .A2(n3611), .ZN(n3645) );
NAND2_X1 U21963 ( .A1(n21366), .A2(n21365), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_27) );
NAND2_X1 U21964 ( .A1(n3642), .A2(n3643), .ZN(n14799) );
NAND2_X1 U21965 ( .A1(n16430), .A2(n15962), .ZN(n3643) );
NAND2_X1 U21966 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_28), .A2(n16429), .ZN(n3642) );
NAND2_X1 U21967 ( .A1(n21370), .A2(n21369), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_28) );
NAND2_X1 U21968 ( .A1(n3639), .A2(n3640), .ZN(n14797) );
NAND2_X1 U21969 ( .A1(n16431), .A2(n15963), .ZN(n3640) );
NAND2_X1 U21970 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_29), .A2(n16429), .ZN(n3639) );
NAND2_X1 U21971 ( .A1(n21373), .A2(n21372), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_29) );
NAND2_X1 U21972 ( .A1(n3633), .A2(n3634), .ZN(n14795) );
NAND2_X1 U21973 ( .A1(n16431), .A2(n15964), .ZN(n3634) );
NAND2_X1 U21974 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_30), .A2(n16429), .ZN(n3633) );
NAND2_X1 U21975 ( .A1(n21379), .A2(n21378), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_30) );
NAND2_X1 U21976 ( .A1(n3630), .A2(n3631), .ZN(n14793) );
NAND2_X1 U21977 ( .A1(n16431), .A2(n15965), .ZN(n3631) );
NAND2_X1 U21978 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_31), .A2(n3611), .ZN(n3630) );
NAND2_X1 U21979 ( .A1(n21383), .A2(n21382), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fetch_addr_d_31) );
NAND2_X1 U21980 ( .A1(n3387), .A2(n3388), .ZN(n15672) );
NAND2_X1 U21981 ( .A1(n3290), .A2(n16124), .ZN(n3388) );
NOR2_X1 U21982 ( .A1(n3390), .A2(n3391), .ZN(n3387) );
NOR2_X1 U21983 ( .A1(n19961), .A2(n3262), .ZN(n3391) );
NAND2_X1 U21984 ( .A1(n3288), .A2(n3289), .ZN(n15670) );
NAND2_X1 U21985 ( .A1(n3290), .A2(n15966), .ZN(n3289) );
NOR2_X1 U21986 ( .A1(n3291), .A2(n3292), .ZN(n3288) );
NOR2_X1 U21987 ( .A1(n19908), .A2(n3262), .ZN(n3292) );
NAND2_X1 U21988 ( .A1(n3293), .A2(n3294), .ZN(n15669) );
NAND2_X1 U21989 ( .A1(n3290), .A2(n15967), .ZN(n3294) );
NOR2_X1 U21990 ( .A1(n3295), .A2(n3296), .ZN(n3293) );
NOR2_X1 U21991 ( .A1(n19911), .A2(n3262), .ZN(n3296) );
NAND2_X1 U21992 ( .A1(n3321), .A2(n3322), .ZN(n15663) );
NAND2_X1 U21993 ( .A1(n3290), .A2(n15968), .ZN(n3322) );
NOR2_X1 U21994 ( .A1(n3323), .A2(n3324), .ZN(n3321) );
NOR2_X1 U21995 ( .A1(n19924), .A2(n16434), .ZN(n3324) );
NAND2_X1 U21996 ( .A1(n3333), .A2(n3334), .ZN(n15660) );
NAND2_X1 U21997 ( .A1(n3290), .A2(n15969), .ZN(n3334) );
NOR2_X1 U21998 ( .A1(n3335), .A2(n3336), .ZN(n3333) );
NOR2_X1 U21999 ( .A1(n19930), .A2(n16434), .ZN(n3336) );
NAND2_X1 U22000 ( .A1(n3353), .A2(n3354), .ZN(n15656) );
NAND2_X1 U22001 ( .A1(n3290), .A2(n16044), .ZN(n3354) );
NOR2_X1 U22002 ( .A1(n3356), .A2(n3357), .ZN(n3353) );
NOR2_X1 U22003 ( .A1(n19944), .A2(n16434), .ZN(n3357) );
NAND2_X1 U22004 ( .A1(n3358), .A2(n3359), .ZN(n15655) );
NAND2_X1 U22005 ( .A1(n3290), .A2(n15970), .ZN(n3359) );
NOR2_X1 U22006 ( .A1(n3361), .A2(n3362), .ZN(n3358) );
NOR2_X1 U22007 ( .A1(n19945), .A2(n16434), .ZN(n3362) );
NAND2_X1 U22008 ( .A1(n3341), .A2(n3342), .ZN(n15625) );
NAND2_X1 U22009 ( .A1(n3290), .A2(n15821), .ZN(n3342) );
NOR2_X1 U22010 ( .A1(n3343), .A2(n3344), .ZN(n3341) );
NOR2_X1 U22011 ( .A1(n19960), .A2(n16434), .ZN(n3344) );
NAND2_X1 U22012 ( .A1(n1588), .A2(n1589), .ZN(n15314) );
NAND2_X1 U22013 ( .A1(n1507), .A2(n15818), .ZN(n1588) );
NAND2_X1 U22014 ( .A1(n1590), .A2(n19963), .ZN(n1589) );
NAND2_X1 U22015 ( .A1(n3027), .A2(n3028), .ZN(n15753) );
NAND2_X1 U22016 ( .A1(n3229), .A2(n3230), .ZN(n15687) );
NAND2_X1 U22017 ( .A1(n3126), .A2(n16117), .ZN(n3230) );
NOR2_X1 U22018 ( .A1(n3231), .A2(n3232), .ZN(n3229) );
NOR2_X1 U22019 ( .A1(n19946), .A2(n3129), .ZN(n3232) );
NAND2_X1 U22020 ( .A1(n3124), .A2(n3125), .ZN(n15681) );
NAND2_X1 U22021 ( .A1(n3126), .A2(n16116), .ZN(n3125) );
NOR2_X1 U22022 ( .A1(n3127), .A2(n3128), .ZN(n3124) );
NOR2_X1 U22023 ( .A1(n19952), .A2(n16436), .ZN(n3128) );
NAND2_X1 U22024 ( .A1(n3131), .A2(n3132), .ZN(n15680) );
NAND2_X1 U22025 ( .A1(n3126), .A2(n15971), .ZN(n3132) );
NOR2_X1 U22026 ( .A1(n3133), .A2(n3134), .ZN(n3131) );
NOR2_X1 U22027 ( .A1(n19953), .A2(n16436), .ZN(n3134) );
NAND2_X1 U22028 ( .A1(n3140), .A2(n3141), .ZN(n15678) );
NAND2_X1 U22029 ( .A1(n3126), .A2(n16045), .ZN(n3141) );
NOR2_X1 U22030 ( .A1(n3142), .A2(n3143), .ZN(n3140) );
NOR2_X1 U22031 ( .A1(n19955), .A2(n16436), .ZN(n3143) );
NAND2_X1 U22032 ( .A1(n3144), .A2(n3145), .ZN(n15677) );
NAND2_X1 U22033 ( .A1(n3126), .A2(n15972), .ZN(n3145) );
NOR2_X1 U22034 ( .A1(n3146), .A2(n3147), .ZN(n3144) );
NOR2_X1 U22035 ( .A1(n19956), .A2(n16436), .ZN(n3147) );
NAND2_X1 U22036 ( .A1(n3152), .A2(n3153), .ZN(n15675) );
NAND2_X1 U22037 ( .A1(n3126), .A2(n16046), .ZN(n3153) );
NOR2_X1 U22038 ( .A1(n3154), .A2(n3155), .ZN(n3152) );
NOR2_X1 U22039 ( .A1(n19958), .A2(n16436), .ZN(n3155) );
NAND2_X1 U22040 ( .A1(n3208), .A2(n3209), .ZN(n15673) );
NAND2_X1 U22041 ( .A1(n3126), .A2(n16118), .ZN(n3209) );
NOR2_X1 U22042 ( .A1(n3210), .A2(n3211), .ZN(n3208) );
NOR2_X1 U22043 ( .A1(n19960), .A2(n3129), .ZN(n3211) );
NAND2_X1 U22044 ( .A1(n2370), .A2(n2371), .ZN(n15579) );
NAND2_X1 U22045 ( .A1(n16455), .A2(n15858), .ZN(n2371) );
NAND2_X1 U22046 ( .A1(n1508), .A2(n1509), .ZN(n15344) );
NAND2_X1 U22047 ( .A1(n1507), .A2(n15822), .ZN(n1508) );
NAND2_X1 U22048 ( .A1(n19963), .A2(alu_adder_result_ex_0), .ZN(n1509) );
NAND2_X1 U22049 ( .A1(n2064), .A2(n2065), .ZN(n15601) );
NAND2_X1 U22050 ( .A1(n16455), .A2(n15804), .ZN(n2065) );
NAND2_X1 U22051 ( .A1(n7835), .A2(n7836), .ZN(n15360) );
NAND2_X1 U22052 ( .A1(n7803), .A2(n15973), .ZN(n7836) );
NAND2_X1 U22053 ( .A1(n16349), .A2(n6896), .ZN(n7835) );
NAND2_X1 U22054 ( .A1(n7801), .A2(n7802), .ZN(n14933) );
NAND2_X1 U22055 ( .A1(n7803), .A2(n15974), .ZN(n7802) );
NAND2_X1 U22056 ( .A1(n16348), .A2(n7185), .ZN(n7801) );
NAND2_X1 U22057 ( .A1(n7846), .A2(n7847), .ZN(n14902) );
NAND2_X1 U22058 ( .A1(n7803), .A2(n15975), .ZN(n7847) );
NAND2_X1 U22059 ( .A1(n16349), .A2(n6943), .ZN(n7846) );
NAND2_X1 U22060 ( .A1(n1584), .A2(n1585), .ZN(n15343) );
NAND2_X1 U22061 ( .A1(data_we_o), .A2(n19963), .ZN(n1585) );
NAND2_X1 U22062 ( .A1(n1507), .A2(n15911), .ZN(n1584) );
NAND2_X1 U22063 ( .A1(n7859), .A2(n7860), .ZN(n15362) );
NAND2_X1 U22064 ( .A1(n7803), .A2(n15976), .ZN(n7860) );
NAND2_X1 U22065 ( .A1(n19977), .A2(n7069), .ZN(n7859) );
NAND2_X1 U22066 ( .A1(n1685), .A2(n1686), .ZN(n15312) );
NAND2_X1 U22067 ( .A1(n16461), .A2(crash_dump_o_32_), .ZN(n1685) );
NAND2_X1 U22068 ( .A1(n1657), .A2(alu_adder_result_ex_0), .ZN(n1686) );
NAND2_X1 U22069 ( .A1(n2365), .A2(n2366), .ZN(n15603) );
NAND2_X1 U22070 ( .A1(n16457), .A2(n15805), .ZN(n2366) );
NAND2_X1 U22071 ( .A1(n8093), .A2(n8094), .ZN(n15561) );
NAND2_X1 U22072 ( .A1(n8083), .A2(n16042), .ZN(n8093) );
NAND2_X1 U22073 ( .A1(n19978), .A2(n7068), .ZN(n8094) );
NAND2_X1 U22074 ( .A1(n7633), .A2(n7634), .ZN(n15764) );
NAND2_X1 U22075 ( .A1(n19975), .A2(n16048), .ZN(n7633) );
NAND2_X1 U22076 ( .A1(n7635), .A2(n7577), .ZN(n7634) );
NAND2_X1 U22077 ( .A1(n7636), .A2(n20874), .ZN(n7635) );
NAND2_X1 U22078 ( .A1(n7608), .A2(n7609), .ZN(n15759) );
NAND2_X1 U22079 ( .A1(n19975), .A2(n16047), .ZN(n7608) );
NAND2_X1 U22080 ( .A1(n7610), .A2(n7577), .ZN(n7609) );
NAND2_X1 U22081 ( .A1(n7611), .A2(n7612), .ZN(n7610) );
NAND2_X1 U22082 ( .A1(n9845), .A2(n9846), .ZN(n15758) );
NAND2_X1 U22083 ( .A1(n9891), .A2(n15926), .ZN(n9845) );
NAND2_X1 U22084 ( .A1(n19970), .A2(n7203), .ZN(n9846) );
NAND2_X1 U22085 ( .A1(n8080), .A2(n8081), .ZN(n15558) );
NAND2_X1 U22086 ( .A1(n8083), .A2(n15909), .ZN(n8080) );
NAND2_X1 U22087 ( .A1(n19978), .A2(n7203), .ZN(n8081) );
NAND2_X1 U22088 ( .A1(n7665), .A2(n7666), .ZN(n15100) );
NAND2_X1 U22089 ( .A1(n19975), .A2(n16049), .ZN(n7665) );
NAND2_X1 U22090 ( .A1(n7667), .A2(n7577), .ZN(n7666) );
NAND2_X1 U22091 ( .A1(n7668), .A2(n7669), .ZN(n7667) );
NAND2_X1 U22092 ( .A1(n7584), .A2(n7585), .ZN(n14936) );
NAND2_X1 U22093 ( .A1(n19975), .A2(n15977), .ZN(n7584) );
NAND2_X1 U22094 ( .A1(n7586), .A2(n7577), .ZN(n7585) );
NAND2_X1 U22095 ( .A1(n7587), .A2(n7588), .ZN(n7586) );
NAND2_X1 U22096 ( .A1(n7592), .A2(n7593), .ZN(n14921) );
NAND2_X1 U22097 ( .A1(n19975), .A2(n16050), .ZN(n7592) );
NAND2_X1 U22098 ( .A1(n7594), .A2(n7577), .ZN(n7593) );
NAND2_X1 U22099 ( .A1(n7595), .A2(n7596), .ZN(n7594) );
NAND2_X1 U22100 ( .A1(n7574), .A2(n7575), .ZN(n14855) );
NAND2_X1 U22101 ( .A1(n19975), .A2(n15978), .ZN(n7574) );
NAND2_X1 U22102 ( .A1(n7576), .A2(n7577), .ZN(n7575) );
NAND2_X1 U22103 ( .A1(n7578), .A2(n7579), .ZN(n7576) );
NAND2_X1 U22104 ( .A1(n2365), .A2(n2676), .ZN(n15602) );
NAND2_X1 U22105 ( .A1(n16456), .A2(n15859), .ZN(n2676) );
NAND2_X1 U22106 ( .A1(n8088), .A2(n8089), .ZN(n15065) );
NAND2_X1 U22107 ( .A1(n8083), .A2(n16043), .ZN(n8088) );
NAND2_X1 U22108 ( .A1(n19978), .A2(n7237), .ZN(n8089) );
NAND2_X1 U22109 ( .A1(n5144), .A2(n5145), .ZN(n15267) );
OR2_X1 U22110 ( .A1(n5146), .A2(n5147), .ZN(n5145) );
NOR2_X1 U22111 ( .A1(n5148), .A2(n5149), .ZN(n5144) );
NOR2_X1 U22112 ( .A1(n19984), .A2(n5151), .ZN(n5149) );
NAND2_X1 U22113 ( .A1(n5106), .A2(n5107), .ZN(n15406) );
NOR2_X1 U22114 ( .A1(n5109), .A2(n5110), .ZN(n5106) );
NOR2_X1 U22115 ( .A1(n15773), .A2(n5108), .ZN(n5107) );
NOR2_X1 U22116 ( .A1(n16125), .A2(n5112), .ZN(n5110) );
NAND2_X1 U22117 ( .A1(n2242), .A2(n2243), .ZN(n15622) );
NAND2_X1 U22118 ( .A1(n16455), .A2(n15820), .ZN(n2243) );
NAND2_X1 U22119 ( .A1(n2412), .A2(n2413), .ZN(n15620) );
NAND2_X1 U22120 ( .A1(n16456), .A2(n15921), .ZN(n2413) );
NAND2_X1 U22121 ( .A1(n2074), .A2(n2075), .ZN(n15616) );
NAND2_X1 U22122 ( .A1(n16455), .A2(n15892), .ZN(n2075) );
NAND2_X1 U22123 ( .A1(n2074), .A2(n2509), .ZN(n15615) );
NAND2_X1 U22124 ( .A1(n16454), .A2(n16128), .ZN(n2509) );
NAND2_X1 U22125 ( .A1(n2084), .A2(n2085), .ZN(n15614) );
NAND2_X1 U22126 ( .A1(n16456), .A2(n15982), .ZN(n2085) );
NAND2_X1 U22127 ( .A1(n2084), .A2(n2558), .ZN(n15613) );
NAND2_X1 U22128 ( .A1(n16455), .A2(n15827), .ZN(n2558) );
NAND2_X1 U22129 ( .A1(n2087), .A2(n2088), .ZN(n15612) );
NAND2_X1 U22130 ( .A1(n16456), .A2(n15815), .ZN(n2088) );
NAND2_X1 U22131 ( .A1(n2087), .A2(n2584), .ZN(n15611) );
NAND2_X1 U22132 ( .A1(n16456), .A2(n15860), .ZN(n2584) );
NAND2_X1 U22133 ( .A1(n2090), .A2(n2091), .ZN(n15610) );
NAND2_X1 U22134 ( .A1(n16455), .A2(n15824), .ZN(n2091) );
NAND2_X1 U22135 ( .A1(n2090), .A2(n2610), .ZN(n15609) );
NAND2_X1 U22136 ( .A1(n16455), .A2(n15914), .ZN(n2610) );
NAND2_X1 U22137 ( .A1(n2064), .A2(n2458), .ZN(n15600) );
NAND2_X1 U22138 ( .A1(n16455), .A2(n15910), .ZN(n2458) );
NAND2_X1 U22139 ( .A1(n2066), .A2(n2067), .ZN(n15599) );
NAND2_X1 U22140 ( .A1(n16457), .A2(n15876), .ZN(n2067) );
NAND2_X1 U22141 ( .A1(n2066), .A2(n2472), .ZN(n15598) );
NAND2_X1 U22142 ( .A1(n16457), .A2(n15908), .ZN(n2472) );
NAND2_X1 U22143 ( .A1(n2093), .A2(n2094), .ZN(n15597) );
NAND2_X1 U22144 ( .A1(n16457), .A2(n15807), .ZN(n2094) );
NAND2_X1 U22145 ( .A1(n2093), .A2(n2640), .ZN(n15596) );
NAND2_X1 U22146 ( .A1(n16456), .A2(n15816), .ZN(n2640) );
NAND2_X1 U22147 ( .A1(n2061), .A2(n2062), .ZN(n15592) );
NAND2_X1 U22148 ( .A1(n16454), .A2(n15917), .ZN(n2062) );
NAND2_X1 U22149 ( .A1(n2061), .A2(n2449), .ZN(n15591) );
NAND2_X1 U22150 ( .A1(n16455), .A2(n15799), .ZN(n2449) );
NAND2_X1 U22151 ( .A1(n2367), .A2(n2368), .ZN(n15588) );
NAND2_X1 U22152 ( .A1(n16454), .A2(n15879), .ZN(n2368) );
NAND2_X1 U22153 ( .A1(n2367), .A2(n2689), .ZN(n15587) );
NAND2_X1 U22154 ( .A1(n16457), .A2(n15810), .ZN(n2689) );
NAND2_X1 U22155 ( .A1(n2068), .A2(n2069), .ZN(n15586) );
NAND2_X1 U22156 ( .A1(n16454), .A2(n15884), .ZN(n2069) );
NAND2_X1 U22157 ( .A1(n2068), .A2(n2489), .ZN(n15585) );
NAND2_X1 U22158 ( .A1(n16456), .A2(n15814), .ZN(n2489) );
NAND2_X1 U22159 ( .A1(n2071), .A2(n2072), .ZN(n15584) );
NAND2_X1 U22160 ( .A1(n16454), .A2(n15924), .ZN(n2072) );
NAND2_X1 U22161 ( .A1(n2071), .A2(n2492), .ZN(n15583) );
NAND2_X1 U22162 ( .A1(n16454), .A2(n16119), .ZN(n2492) );
NAND2_X1 U22163 ( .A1(n2081), .A2(n2082), .ZN(n15582) );
NAND2_X1 U22164 ( .A1(n16455), .A2(n15918), .ZN(n2082) );
NAND2_X1 U22165 ( .A1(n2370), .A2(n2705), .ZN(n15578) );
NAND2_X1 U22166 ( .A1(n16457), .A2(n15893), .ZN(n2705) );
NAND2_X1 U22167 ( .A1(n9892), .A2(n9893), .ZN(n15756) );
NAND2_X1 U22168 ( .A1(n9891), .A2(n15979), .ZN(n9892) );
NAND2_X1 U22169 ( .A1(n19970), .A2(n7253), .ZN(n9893) );
NAND2_X1 U22170 ( .A1(n2245), .A2(n2246), .ZN(n15580) );
NOR2_X1 U22171 ( .A1(n2258), .A2(n2259), .ZN(n2245) );
NOR2_X1 U22172 ( .A1(n19877), .A2(n2248), .ZN(n2246) );
AND2_X1 U22173 ( .A1(n2103), .A2(n2261), .ZN(n2258) );
NAND2_X1 U22174 ( .A1(n5573), .A2(n5574), .ZN(n15554) );
NAND2_X1 U22175 ( .A1(n5571), .A2(n15823), .ZN(n5573) );
NAND2_X1 U22176 ( .A1(n20911), .A2(n5575), .ZN(n5574) );
NAND2_X1 U22177 ( .A1(n15811), .A2(n5087), .ZN(n5575) );
NAND2_X1 U22178 ( .A1(n5566), .A2(n5567), .ZN(n15553) );
NAND2_X1 U22179 ( .A1(n5571), .A2(n15922), .ZN(n5566) );
NAND2_X1 U22180 ( .A1(n20911), .A2(n5569), .ZN(n5567) );
NAND2_X1 U22181 ( .A1(n15811), .A2(n4959), .ZN(n5569) );
NAND2_X1 U22182 ( .A1(n1532), .A2(n1533), .ZN(n15551) );
NAND2_X1 U22183 ( .A1(n1534), .A2(n15825), .ZN(n1533) );
NOR2_X1 U22184 ( .A1(n1538), .A2(n1539), .ZN(n1532) );
NAND2_X1 U22185 ( .A1(n1531), .A2(n1536), .ZN(n1534) );
NAND2_X1 U22186 ( .A1(n4942), .A2(n4943), .ZN(n15419) );
NOR2_X1 U22187 ( .A1(n5083), .A2(n5084), .ZN(n4942) );
NOR2_X1 U22188 ( .A1(n4944), .A2(n4945), .ZN(n4943) );
NOR2_X1 U22189 ( .A1(n20681), .A2(n4936), .ZN(n5084) );
NAND2_X1 U22190 ( .A1(n2217), .A2(n2218), .ZN(n15606) );
NOR2_X1 U22191 ( .A1(n2239), .A2(n2240), .ZN(n2217) );
NOR2_X1 U22192 ( .A1(n2219), .A2(n2220), .ZN(n2218) );
NOR2_X1 U22193 ( .A1(n16457), .A2(n2241), .ZN(n2239) );
NAND2_X1 U22194 ( .A1(n1555), .A2(n1556), .ZN(n15547) );
NAND2_X1 U22195 ( .A1(n1567), .A2(n15916), .ZN(n1555) );
NAND2_X1 U22196 ( .A1(n19964), .A2(n1558), .ZN(n1556) );
INV_X1 U22197 ( .A(n1567), .ZN(n19964) );
NAND2_X1 U22198 ( .A1(n5174), .A2(n5175), .ZN(n15560) );
NOR2_X1 U22199 ( .A1(n5183), .A2(n5184), .ZN(n5174) );
NOR2_X1 U22200 ( .A1(n5176), .A2(n5177), .ZN(n5175) );
NAND2_X1 U22201 ( .A1(n5178), .A2(n20873), .ZN(n5177) );
NAND2_X1 U22202 ( .A1(n2130), .A2(n2131), .ZN(n15608) );
NOR2_X1 U22203 ( .A1(n2154), .A2(n2155), .ZN(n2130) );
NOR2_X1 U22204 ( .A1(n2132), .A2(n2133), .ZN(n2131) );
NAND2_X1 U22205 ( .A1(n2156), .A2(n2157), .ZN(n2155) );
NAND2_X1 U22206 ( .A1(n6752), .A2(n6753), .ZN(n15262) );
AND2_X1 U22207 ( .A1(n6754), .A2(n6755), .ZN(n6753) );
NOR2_X1 U22208 ( .A1(n6759), .A2(n6760), .ZN(n6752) );
NAND2_X1 U22209 ( .A1(id_stage_i_controller_i_N262), .A2(n16403), .ZN(n6755) );
NAND2_X1 U22210 ( .A1(n6774), .A2(n6775), .ZN(n15261) );
AND2_X1 U22211 ( .A1(n6776), .A2(n6777), .ZN(n6775) );
NOR2_X1 U22212 ( .A1(n6781), .A2(n6782), .ZN(n6774) );
NAND2_X1 U22213 ( .A1(id_stage_i_controller_i_N260), .A2(n16403), .ZN(n6777) );
NAND2_X1 U22214 ( .A1(n6704), .A2(n6705), .ZN(n14984) );
AND2_X1 U22215 ( .A1(n6706), .A2(n6707), .ZN(n6705) );
NOR2_X1 U22216 ( .A1(n6713), .A2(n6714), .ZN(n6704) );
NAND2_X1 U22217 ( .A1(id_stage_i_controller_i_N266), .A2(n16403), .ZN(n6707) );
NAND2_X1 U22218 ( .A1(n6720), .A2(n6721), .ZN(n14970) );
AND2_X1 U22219 ( .A1(n6722), .A2(n6723), .ZN(n6721) );
NOR2_X1 U22220 ( .A1(n6726), .A2(n6727), .ZN(n6720) );
NAND2_X1 U22221 ( .A1(id_stage_i_controller_i_N265), .A2(n16403), .ZN(n6723) );
NAND2_X1 U22222 ( .A1(n6741), .A2(n6742), .ZN(n14956) );
AND2_X1 U22223 ( .A1(n6743), .A2(n6744), .ZN(n6742) );
NOR2_X1 U22224 ( .A1(n6748), .A2(n6749), .ZN(n6741) );
NAND2_X1 U22225 ( .A1(id_stage_i_controller_i_N263), .A2(n16403), .ZN(n6744) );
NAND2_X1 U22226 ( .A1(n6763), .A2(n6764), .ZN(n14943) );
AND2_X1 U22227 ( .A1(n6765), .A2(n6766), .ZN(n6764) );
NOR2_X1 U22228 ( .A1(n6770), .A2(n6771), .ZN(n6763) );
NAND2_X1 U22229 ( .A1(id_stage_i_controller_i_N261), .A2(n16403), .ZN(n6766) );
NAND2_X1 U22230 ( .A1(n6730), .A2(n6731), .ZN(n14931) );
AND2_X1 U22231 ( .A1(n6732), .A2(n6733), .ZN(n6731) );
NOR2_X1 U22232 ( .A1(n6737), .A2(n6738), .ZN(n6730) );
NAND2_X1 U22233 ( .A1(id_stage_i_controller_i_N264), .A2(n16403), .ZN(n6733) );
NAND2_X1 U22234 ( .A1(n6806), .A2(n6807), .ZN(n15260) );
AND2_X1 U22235 ( .A1(n6808), .A2(n6809), .ZN(n6807) );
NOR2_X1 U22236 ( .A1(n6813), .A2(n6814), .ZN(n6806) );
NAND2_X1 U22237 ( .A1(id_stage_i_controller_i_N259), .A2(n6708), .ZN(n6809) );
NAND2_X1 U22238 ( .A1(n6908), .A2(n6909), .ZN(n15258) );
AND2_X1 U22239 ( .A1(n6910), .A2(n6911), .ZN(n6909) );
NOR2_X1 U22240 ( .A1(n6915), .A2(n6916), .ZN(n6908) );
NAND2_X1 U22241 ( .A1(id_stage_i_controller_i_N258), .A2(n6708), .ZN(n6911) );
NAND2_X1 U22242 ( .A1(n6985), .A2(n6986), .ZN(n15257) );
AND2_X1 U22243 ( .A1(n6987), .A2(n6988), .ZN(n6986) );
NOR2_X1 U22244 ( .A1(n6991), .A2(n6992), .ZN(n6985) );
NAND2_X1 U22245 ( .A1(id_stage_i_controller_i_N269), .A2(n6708), .ZN(n6988) );
NAND2_X1 U22246 ( .A1(n6995), .A2(n6996), .ZN(n15256) );
AND2_X1 U22247 ( .A1(n6997), .A2(n6998), .ZN(n6996) );
NOR2_X1 U22248 ( .A1(n7001), .A2(n7002), .ZN(n6995) );
NAND2_X1 U22249 ( .A1(id_stage_i_controller_i_N268), .A2(n6708), .ZN(n6998) );
NAND2_X1 U22250 ( .A1(n6955), .A2(n6956), .ZN(n15066) );
AND2_X1 U22251 ( .A1(n6957), .A2(n6958), .ZN(n6956) );
NOR2_X1 U22252 ( .A1(n6961), .A2(n6962), .ZN(n6955) );
NAND2_X1 U22253 ( .A1(id_stage_i_controller_i_N272), .A2(n16403), .ZN(n6958) );
NAND2_X1 U22254 ( .A1(n6965), .A2(n6966), .ZN(n15051) );
AND2_X1 U22255 ( .A1(n6967), .A2(n6968), .ZN(n6966) );
NOR2_X1 U22256 ( .A1(n6971), .A2(n6972), .ZN(n6965) );
NAND2_X1 U22257 ( .A1(id_stage_i_controller_i_N271), .A2(n6708), .ZN(n6968) );
NAND2_X1 U22258 ( .A1(n6975), .A2(n6976), .ZN(n15037) );
AND2_X1 U22259 ( .A1(n6977), .A2(n6978), .ZN(n6976) );
NOR2_X1 U22260 ( .A1(n6981), .A2(n6982), .ZN(n6975) );
NAND2_X1 U22261 ( .A1(id_stage_i_controller_i_N270), .A2(n16403), .ZN(n6978) );
NAND2_X1 U22262 ( .A1(n7005), .A2(n7006), .ZN(n14998) );
AND2_X1 U22263 ( .A1(n7007), .A2(n7008), .ZN(n7006) );
NOR2_X1 U22264 ( .A1(n7011), .A2(n7012), .ZN(n7005) );
NAND2_X1 U22265 ( .A1(id_stage_i_controller_i_N267), .A2(n6708), .ZN(n7008) );
NAND2_X1 U22266 ( .A1(n4749), .A2(n4750), .ZN(n15434) );
NOR2_X1 U22267 ( .A1(n4760), .A2(n4761), .ZN(n4749) );
NOR2_X1 U22268 ( .A1(n4751), .A2(n4752), .ZN(n4750) );
NAND2_X1 U22269 ( .A1(n4762), .A2(n4763), .ZN(n4761) );
NAND2_X1 U22270 ( .A1(n4689), .A2(n4690), .ZN(n15432) );
NOR2_X1 U22271 ( .A1(n4700), .A2(n4701), .ZN(n4689) );
NOR2_X1 U22272 ( .A1(n4691), .A2(n4692), .ZN(n4690) );
NAND2_X1 U22273 ( .A1(n4702), .A2(n4703), .ZN(n4701) );
NAND2_X1 U22274 ( .A1(n4668), .A2(n4669), .ZN(n15431) );
NOR2_X1 U22275 ( .A1(n4679), .A2(n4680), .ZN(n4668) );
NOR2_X1 U22276 ( .A1(n4670), .A2(n4671), .ZN(n4669) );
NAND2_X1 U22277 ( .A1(n4681), .A2(n4682), .ZN(n4680) );
NAND2_X1 U22278 ( .A1(n4626), .A2(n4627), .ZN(n15429) );
NOR2_X1 U22279 ( .A1(n4637), .A2(n4638), .ZN(n4626) );
NOR2_X1 U22280 ( .A1(n4628), .A2(n4629), .ZN(n4627) );
NAND2_X1 U22281 ( .A1(n4639), .A2(n4640), .ZN(n4638) );
NAND2_X1 U22282 ( .A1(n4436), .A2(n4437), .ZN(n15471) );
NOR2_X1 U22283 ( .A1(n4450), .A2(n4451), .ZN(n4436) );
NOR2_X1 U22284 ( .A1(n4438), .A2(n4439), .ZN(n4437) );
NAND2_X1 U22285 ( .A1(n4452), .A2(n4453), .ZN(n4451) );
NAND2_X1 U22286 ( .A1(n4791), .A2(n4792), .ZN(n15436) );
NOR2_X1 U22287 ( .A1(n4803), .A2(n4804), .ZN(n4791) );
NOR2_X1 U22288 ( .A1(n4793), .A2(n4794), .ZN(n4792) );
NAND2_X1 U22289 ( .A1(n4805), .A2(n4806), .ZN(n4804) );
NAND2_X1 U22290 ( .A1(n4770), .A2(n4771), .ZN(n15435) );
NOR2_X1 U22291 ( .A1(n4781), .A2(n4782), .ZN(n4770) );
NOR2_X1 U22292 ( .A1(n4772), .A2(n4773), .ZN(n4771) );
NAND2_X1 U22293 ( .A1(n4783), .A2(n4784), .ZN(n4782) );
NAND2_X1 U22294 ( .A1(n4728), .A2(n4729), .ZN(n15433) );
NOR2_X1 U22295 ( .A1(n4739), .A2(n4740), .ZN(n4728) );
NOR2_X1 U22296 ( .A1(n4730), .A2(n4731), .ZN(n4729) );
NAND2_X1 U22297 ( .A1(n4741), .A2(n4742), .ZN(n4740) );
NAND2_X1 U22298 ( .A1(n4647), .A2(n4648), .ZN(n15430) );
NOR2_X1 U22299 ( .A1(n4658), .A2(n4659), .ZN(n4647) );
NOR2_X1 U22300 ( .A1(n4649), .A2(n4650), .ZN(n4648) );
NAND2_X1 U22301 ( .A1(n4660), .A2(n4661), .ZN(n4659) );
NAND2_X1 U22302 ( .A1(n4605), .A2(n4606), .ZN(n15428) );
NOR2_X1 U22303 ( .A1(n4616), .A2(n4617), .ZN(n4605) );
NOR2_X1 U22304 ( .A1(n4607), .A2(n4608), .ZN(n4606) );
NAND2_X1 U22305 ( .A1(n4618), .A2(n4619), .ZN(n4617) );
NAND2_X1 U22306 ( .A1(n4584), .A2(n4585), .ZN(n15427) );
NOR2_X1 U22307 ( .A1(n4595), .A2(n4596), .ZN(n4584) );
NOR2_X1 U22308 ( .A1(n4586), .A2(n4587), .ZN(n4585) );
NAND2_X1 U22309 ( .A1(n4597), .A2(n4598), .ZN(n4596) );
NAND2_X1 U22310 ( .A1(n4563), .A2(n4564), .ZN(n15426) );
NOR2_X1 U22311 ( .A1(n4574), .A2(n4575), .ZN(n4563) );
NOR2_X1 U22312 ( .A1(n4565), .A2(n4566), .ZN(n4564) );
NAND2_X1 U22313 ( .A1(n4576), .A2(n4577), .ZN(n4575) );
NAND2_X1 U22314 ( .A1(n4542), .A2(n4543), .ZN(n15425) );
NOR2_X1 U22315 ( .A1(n4553), .A2(n4554), .ZN(n4542) );
NOR2_X1 U22316 ( .A1(n4544), .A2(n4545), .ZN(n4543) );
NAND2_X1 U22317 ( .A1(n4555), .A2(n4556), .ZN(n4554) );
NAND2_X1 U22318 ( .A1(n4521), .A2(n4522), .ZN(n15424) );
NOR2_X1 U22319 ( .A1(n4532), .A2(n4533), .ZN(n4521) );
NOR2_X1 U22320 ( .A1(n4523), .A2(n4524), .ZN(n4522) );
NAND2_X1 U22321 ( .A1(n4534), .A2(n4535), .ZN(n4533) );
NAND2_X1 U22322 ( .A1(n4500), .A2(n4501), .ZN(n15423) );
NOR2_X1 U22323 ( .A1(n4511), .A2(n4512), .ZN(n4500) );
NOR2_X1 U22324 ( .A1(n4502), .A2(n4503), .ZN(n4501) );
NAND2_X1 U22325 ( .A1(n4513), .A2(n4514), .ZN(n4512) );
NAND2_X1 U22326 ( .A1(n4460), .A2(n4461), .ZN(n15422) );
NOR2_X1 U22327 ( .A1(n4471), .A2(n4472), .ZN(n4460) );
NOR2_X1 U22328 ( .A1(n4462), .A2(n4463), .ZN(n4461) );
NAND2_X1 U22329 ( .A1(n4473), .A2(n4474), .ZN(n4472) );
NAND2_X1 U22330 ( .A1(n4870), .A2(n4871), .ZN(n15440) );
NOR2_X1 U22331 ( .A1(n4879), .A2(n4880), .ZN(n4870) );
NOR2_X1 U22332 ( .A1(n4872), .A2(n4873), .ZN(n4871) );
NAND2_X1 U22333 ( .A1(n4881), .A2(n4882), .ZN(n4880) );
NAND2_X1 U22334 ( .A1(n4851), .A2(n4852), .ZN(n15439) );
NOR2_X1 U22335 ( .A1(n4860), .A2(n4861), .ZN(n4851) );
NOR2_X1 U22336 ( .A1(n4853), .A2(n4854), .ZN(n4852) );
NAND2_X1 U22337 ( .A1(n4862), .A2(n4863), .ZN(n4861) );
NAND2_X1 U22338 ( .A1(n4832), .A2(n4833), .ZN(n15438) );
NOR2_X1 U22339 ( .A1(n4841), .A2(n4842), .ZN(n4832) );
NOR2_X1 U22340 ( .A1(n4834), .A2(n4835), .ZN(n4833) );
NAND2_X1 U22341 ( .A1(n4843), .A2(n4844), .ZN(n4842) );
NAND2_X1 U22342 ( .A1(n4813), .A2(n4814), .ZN(n15437) );
NOR2_X1 U22343 ( .A1(n4822), .A2(n4823), .ZN(n4813) );
NOR2_X1 U22344 ( .A1(n4815), .A2(n4816), .ZN(n4814) );
NAND2_X1 U22345 ( .A1(n4824), .A2(n4825), .ZN(n4823) );
NAND2_X1 U22346 ( .A1(n4908), .A2(n4909), .ZN(n15472) );
NOR2_X1 U22347 ( .A1(n4920), .A2(n4921), .ZN(n4908) );
NOR2_X1 U22348 ( .A1(n4910), .A2(n4911), .ZN(n4909) );
NAND2_X1 U22349 ( .A1(n4922), .A2(n4923), .ZN(n4921) );
NAND2_X1 U22350 ( .A1(n4889), .A2(n4890), .ZN(n15441) );
NOR2_X1 U22351 ( .A1(n4898), .A2(n4899), .ZN(n4889) );
NOR2_X1 U22352 ( .A1(n4891), .A2(n4892), .ZN(n4890) );
NAND2_X1 U22353 ( .A1(n4900), .A2(n4901), .ZN(n4899) );
NAND2_X1 U22354 ( .A1(n4710), .A2(n4711), .ZN(n15418) );
NOR2_X1 U22355 ( .A1(n4719), .A2(n4720), .ZN(n4710) );
NOR2_X1 U22356 ( .A1(n4712), .A2(n4713), .ZN(n4711) );
NAND2_X1 U22357 ( .A1(n4721), .A2(n4722), .ZN(n4720) );
NAND2_X1 U22358 ( .A1(n4481), .A2(n4482), .ZN(n15417) );
NOR2_X1 U22359 ( .A1(n4490), .A2(n4491), .ZN(n4481) );
NOR2_X1 U22360 ( .A1(n4483), .A2(n4484), .ZN(n4482) );
NAND2_X1 U22361 ( .A1(n4492), .A2(n4493), .ZN(n4491) );
NAND2_X1 U22362 ( .A1(n4387), .A2(n4388), .ZN(n15416) );
NOR2_X1 U22363 ( .A1(n4396), .A2(n4397), .ZN(n4387) );
NOR2_X1 U22364 ( .A1(n4389), .A2(n4390), .ZN(n4388) );
NAND2_X1 U22365 ( .A1(n4398), .A2(n4399), .ZN(n4397) );
NAND2_X1 U22366 ( .A1(n4368), .A2(n4369), .ZN(n15415) );
NOR2_X1 U22367 ( .A1(n4377), .A2(n4378), .ZN(n4368) );
NOR2_X1 U22368 ( .A1(n4370), .A2(n4371), .ZN(n4369) );
NAND2_X1 U22369 ( .A1(n4379), .A2(n4380), .ZN(n4378) );
NAND2_X1 U22370 ( .A1(n4349), .A2(n4350), .ZN(n15414) );
NOR2_X1 U22371 ( .A1(n4358), .A2(n4359), .ZN(n4349) );
NOR2_X1 U22372 ( .A1(n4351), .A2(n4352), .ZN(n4350) );
NAND2_X1 U22373 ( .A1(n4360), .A2(n4361), .ZN(n4359) );
NAND2_X1 U22374 ( .A1(n4330), .A2(n4331), .ZN(n15413) );
NOR2_X1 U22375 ( .A1(n4339), .A2(n4340), .ZN(n4330) );
NOR2_X1 U22376 ( .A1(n4332), .A2(n4333), .ZN(n4331) );
NAND2_X1 U22377 ( .A1(n4341), .A2(n4342), .ZN(n4340) );
NAND2_X1 U22378 ( .A1(n4311), .A2(n4312), .ZN(n15412) );
NOR2_X1 U22379 ( .A1(n4320), .A2(n4321), .ZN(n4311) );
NOR2_X1 U22380 ( .A1(n4313), .A2(n4314), .ZN(n4312) );
NAND2_X1 U22381 ( .A1(n4322), .A2(n4323), .ZN(n4321) );
NAND2_X1 U22382 ( .A1(n4292), .A2(n4293), .ZN(n15411) );
NOR2_X1 U22383 ( .A1(n4301), .A2(n4302), .ZN(n4292) );
NOR2_X1 U22384 ( .A1(n4294), .A2(n4295), .ZN(n4293) );
NAND2_X1 U22385 ( .A1(n4303), .A2(n4304), .ZN(n4302) );
NAND2_X1 U22386 ( .A1(n4262), .A2(n4263), .ZN(n15410) );
NOR2_X1 U22387 ( .A1(n4276), .A2(n4277), .ZN(n4262) );
NOR2_X1 U22388 ( .A1(n4264), .A2(n4265), .ZN(n4263) );
NAND2_X1 U22389 ( .A1(n4278), .A2(n4279), .ZN(n4277) );
NAND2_X1 U22390 ( .A1(n3045), .A2(n19882), .ZN(n15741) );
INV_X1 U22391 ( .A(n3036), .ZN(n19882) );
NOR2_X1 U22392 ( .A1(n3052), .A2(n3053), .ZN(n3045) );
AND2_X1 U22393 ( .A1(n3041), .A2(n19885), .ZN(n3053) );
AND2_X1 U22394 ( .A1(n16130), .A2(n1511), .ZN(n15550) );
NAND2_X1 U22395 ( .A1(rf_rdata_b_ecc_i_15_), .A2(n5586), .ZN(n5604) );
NAND2_X1 U22396 ( .A1(rf_rdata_b_ecc_i_31_), .A2(n5272), .ZN(n5603) );
OR2_X4 U22397 ( .A1(n16268), .A2(n16269), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0) );
AND2_X1 U22398 ( .A1(rf_rdata_a_ecc_i_16_), .A2(n5274), .ZN(n16268) );
AND2_X1 U22399 ( .A1(rf_rdata_a_ecc_i_0_), .A2(n11299), .ZN(n16269) );
NAND2_X1 U22400 ( .A1(rf_rdata_b_ecc_i_17_), .A2(n5272), .ZN(n5601) );
NAND2_X1 U22401 ( .A1(rf_rdata_b_ecc_i_1_), .A2(n5586), .ZN(n5602) );
NAND2_X2 U22402 ( .A1(n5629), .A2(n5630), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3) );
NAND2_X1 U22403 ( .A1(rf_rdata_a_ecc_i_3_), .A2(n11299), .ZN(n5629) );
NAND2_X1 U22404 ( .A1(rf_rdata_a_ecc_i_19_), .A2(n5274), .ZN(n5630) );
NAND2_X2 U22405 ( .A1(n5627), .A2(n5628), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4) );
NAND2_X1 U22406 ( .A1(rf_rdata_a_ecc_i_4_), .A2(n11299), .ZN(n5627) );
NAND2_X1 U22407 ( .A1(rf_rdata_a_ecc_i_20_), .A2(n5274), .ZN(n5628) );
NAND2_X2 U22408 ( .A1(n5625), .A2(n5626), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5) );
NAND2_X1 U22409 ( .A1(rf_rdata_a_ecc_i_5_), .A2(n11299), .ZN(n5625) );
NAND2_X1 U22410 ( .A1(rf_rdata_a_ecc_i_21_), .A2(n5274), .ZN(n5626) );
NAND2_X2 U22411 ( .A1(n5605), .A2(n5606), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14) );
NAND2_X1 U22412 ( .A1(rf_rdata_b_ecc_i_30_), .A2(n5272), .ZN(n5605) );
NAND2_X1 U22413 ( .A1(rf_rdata_b_ecc_i_14_), .A2(n5586), .ZN(n5606) );
NAND2_X1 U22414 ( .A1(rf_rdata_b_ecc_i_18_), .A2(n5272), .ZN(n5599) );
NAND2_X1 U22415 ( .A1(rf_rdata_b_ecc_i_2_), .A2(n5586), .ZN(n5600) );
NAND2_X1 U22416 ( .A1(rf_rdata_b_ecc_i_19_), .A2(n5272), .ZN(n5597) );
NAND2_X1 U22417 ( .A1(rf_rdata_b_ecc_i_3_), .A2(n5586), .ZN(n5598) );
NAND2_X1 U22418 ( .A1(rf_rdata_b_ecc_i_20_), .A2(n5272), .ZN(n5595) );
NAND2_X1 U22419 ( .A1(rf_rdata_b_ecc_i_4_), .A2(n5586), .ZN(n5596) );
NAND2_X1 U22420 ( .A1(rf_rdata_b_ecc_i_21_), .A2(n5272), .ZN(n5593) );
NAND2_X1 U22421 ( .A1(rf_rdata_b_ecc_i_5_), .A2(n5586), .ZN(n5594) );
NAND2_X1 U22422 ( .A1(rf_rdata_b_ecc_i_22_), .A2(n5272), .ZN(n5591) );
NAND2_X1 U22423 ( .A1(rf_rdata_b_ecc_i_6_), .A2(n5586), .ZN(n5592) );
NAND2_X1 U22424 ( .A1(rf_rdata_b_ecc_i_23_), .A2(n5272), .ZN(n5589) );
NAND2_X1 U22425 ( .A1(rf_rdata_b_ecc_i_7_), .A2(n5586), .ZN(n5590) );
NAND2_X1 U22426 ( .A1(rf_rdata_b_ecc_i_24_), .A2(n5272), .ZN(n5587) );
NAND2_X1 U22427 ( .A1(rf_rdata_b_ecc_i_8_), .A2(n5586), .ZN(n5588) );
NAND2_X1 U22428 ( .A1(rf_rdata_b_ecc_i_25_), .A2(n5272), .ZN(n5584) );
NAND2_X1 U22429 ( .A1(rf_rdata_b_ecc_i_9_), .A2(n5586), .ZN(n5585) );
NAND2_X1 U22430 ( .A1(rf_rdata_b_ecc_i_26_), .A2(n5272), .ZN(n5613) );
NAND2_X1 U22431 ( .A1(rf_rdata_b_ecc_i_10_), .A2(n5586), .ZN(n5614) );
NAND2_X1 U22432 ( .A1(rf_rdata_b_ecc_i_27_), .A2(n5272), .ZN(n5611) );
NAND2_X1 U22433 ( .A1(rf_rdata_b_ecc_i_11_), .A2(n5586), .ZN(n5612) );
NAND2_X1 U22434 ( .A1(rf_rdata_b_ecc_i_28_), .A2(n5272), .ZN(n5609) );
NAND2_X1 U22435 ( .A1(rf_rdata_b_ecc_i_12_), .A2(n5586), .ZN(n5610) );
NAND2_X2 U22436 ( .A1(n5607), .A2(n5608), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13) );
NAND2_X1 U22437 ( .A1(rf_rdata_b_ecc_i_29_), .A2(n5272), .ZN(n5607) );
NAND2_X1 U22438 ( .A1(rf_rdata_b_ecc_i_13_), .A2(n5586), .ZN(n5608) );
NAND2_X1 U22439 ( .A1(rf_rdata_a_ecc_i_2_), .A2(n11299), .ZN(n5631) );
NAND2_X1 U22440 ( .A1(rf_rdata_a_ecc_i_18_), .A2(n5274), .ZN(n5632) );
NAND2_X2 U22441 ( .A1(n5615), .A2(n5616), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0) );
NAND2_X1 U22442 ( .A1(rf_rdata_b_ecc_i_16_), .A2(n5272), .ZN(n5615) );
NAND2_X1 U22443 ( .A1(rf_rdata_b_ecc_i_0_), .A2(n5586), .ZN(n5616) );
NAND2_X1 U22444 ( .A1(n9959), .A2(n9960), .ZN(n1391) );
NOR2_X1 U22445 ( .A1(n9963), .A2(n9964), .ZN(n9959) );
NOR2_X1 U22446 ( .A1(n11061), .A2(n8600), .ZN(n9964) );
NAND2_X1 U22447 ( .A1(n10496), .A2(n10051), .ZN(n10495) );
NAND2_X1 U22448 ( .A1(rf_rdata_b_ecc_i_1_), .A2(n20950), .ZN(n10494) );
NAND2_X1 U22449 ( .A1(n10497), .A2(n10498), .ZN(n10496) );
NAND2_X1 U22450 ( .A1(n10483), .A2(n10484), .ZN(alu_operand_b_ex_2) );
NAND2_X1 U22451 ( .A1(n10485), .A2(n10051), .ZN(n10484) );
NAND2_X1 U22452 ( .A1(rf_rdata_b_ecc_i_2_), .A2(n20950), .ZN(n10483) );
NAND2_X1 U22453 ( .A1(n10486), .A2(n10487), .ZN(n10485) );
NAND2_X1 U22454 ( .A1(n10477), .A2(n10478), .ZN(alu_operand_b_ex_3) );
NOR2_X1 U22455 ( .A1(n10479), .A2(n10480), .ZN(n10477) );
NAND2_X1 U22456 ( .A1(rf_rdata_b_ecc_i_3_), .A2(n16356), .ZN(n10478) );
NOR2_X1 U22457 ( .A1(n11332), .A2(n10158), .ZN(n10479) );
NAND2_X1 U22458 ( .A1(n10507), .A2(n10508), .ZN(ex_block_i_alu_i_shift_amt_compl_0) );
NAND2_X1 U22459 ( .A1(n10509), .A2(n10051), .ZN(n10508) );
NAND2_X1 U22460 ( .A1(rf_rdata_b_ecc_i_0_), .A2(n20950), .ZN(n10507) );
NAND2_X1 U22461 ( .A1(n10510), .A2(n10511), .ZN(n10509) );
NAND2_X1 U22462 ( .A1(n9885), .A2(n9886), .ZN(n466) );
NOR2_X1 U22463 ( .A1(n9889), .A2(n9890), .ZN(n9885) );
NOR2_X1 U22464 ( .A1(n9887), .A2(n9888), .ZN(n9886) );
NOR2_X1 U22465 ( .A1(n11032), .A2(n8600), .ZN(n9890) );
INV_X1 U22466 ( .A(rf_rdata_b_ecc_i_31_), .ZN(n20764) );
INV_X1 U22467 ( .A(n23779), .ZN(n20167) );
INV_X1 U22468 ( .A(n22928), .ZN(n20553) );
INV_X1 U22469 ( .A(n23128), .ZN(n20549) );
INV_X1 U22470 ( .A(n23239), .ZN(n20467) );
INV_X1 U22471 ( .A(n23346), .ZN(n20316) );
INV_X1 U22472 ( .A(n23362), .ZN(n20390) );
INV_X1 U22473 ( .A(n23496), .ZN(n20314) );
INV_X1 U22474 ( .A(n23635), .ZN(n20239) );
INV_X1 U22475 ( .A(n23799), .ZN(n20237) );
INV_X1 U22476 ( .A(rf_rdata_a_ecc_i_0_), .ZN(n20760) );
INV_X1 U22477 ( .A(rf_rdata_a_ecc_i_2_), .ZN(n20752) );
INV_X1 U22478 ( .A(rf_rdata_a_ecc_i_4_), .ZN(n20741) );
INV_X1 U22479 ( .A(rf_rdata_a_ecc_i_3_), .ZN(n20746) );
INV_X1 U22480 ( .A(rf_rdata_a_ecc_i_1_), .ZN(n20756) );
NAND2_X1 U22481 ( .A1(rf_rdata_a_ecc_i_1_), .A2(n11299), .ZN(n5633) );
NAND2_X1 U22482 ( .A1(rf_rdata_a_ecc_i_17_), .A2(n5274), .ZN(n5634) );
NAND2_X1 U22483 ( .A1(n5866), .A2(n5867), .ZN(n5865) );
NAND2_X1 U22484 ( .A1(n11246), .A2(n20960), .ZN(n5867) );
NAND2_X1 U22485 ( .A1(n16409), .A2(n20853), .ZN(n5866) );
NAND2_X1 U22486 ( .A1(n6084), .A2(n6085), .ZN(ex_block_i_alu_i_adder_in_b_1) );
NOR2_X1 U22487 ( .A1(n6086), .A2(n6087), .ZN(n6085) );
NOR2_X1 U22488 ( .A1(n6090), .A2(n6091), .ZN(n6084) );
NOR2_X1 U22489 ( .A1(rf_rdata_b_ecc_i_0_), .A2(n20959), .ZN(n6086) );
NAND2_X1 U22490 ( .A1(n5868), .A2(n5869), .ZN(ex_block_i_alu_i_adder_in_b_4) );
NOR2_X1 U22491 ( .A1(n5870), .A2(n5871), .ZN(n5869) );
NOR2_X1 U22492 ( .A1(n5874), .A2(n5875), .ZN(n5868) );
NOR2_X1 U22493 ( .A1(rf_rdata_b_ecc_i_3_), .A2(n20959), .ZN(n5870) );
INV_X1 U22494 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N36), .ZN(n20673) );
INV_X1 U22495 ( .A(n22860), .ZN(n20552) );
INV_X1 U22496 ( .A(n22870), .ZN(n20590) );
INV_X1 U22497 ( .A(n24045), .ZN(n20572) );
INV_X1 U22498 ( .A(n23044), .ZN(n20586) );
INV_X1 U22499 ( .A(n22567), .ZN(n20602) );
INV_X1 U22500 ( .A(n22645), .ZN(n20562) );
INV_X1 U22501 ( .A(n22654), .ZN(n20600) );
INV_X1 U22502 ( .A(n22614), .ZN(n20560) );
INV_X1 U22503 ( .A(n22624), .ZN(n20598) );
INV_X1 U22504 ( .A(n22768), .ZN(n20558) );
INV_X1 U22505 ( .A(n22777), .ZN(n20596) );
INV_X1 U22506 ( .A(n22715), .ZN(n20556) );
INV_X1 U22507 ( .A(n22725), .ZN(n20594) );
INV_X1 U22508 ( .A(n22929), .ZN(n20516) );
INV_X1 U22509 ( .A(n22936), .ZN(n20554) );
INV_X1 U22510 ( .A(n22945), .ZN(n20592) );
INV_X1 U22511 ( .A(n23129), .ZN(n20512) );
INV_X1 U22512 ( .A(n23136), .ZN(n20550) );
INV_X1 U22513 ( .A(n23145), .ZN(n20588) );
INV_X1 U22514 ( .A(n23256), .ZN(n20506) );
INV_X1 U22515 ( .A(n23263), .ZN(n20544) );
INV_X1 U22516 ( .A(n23272), .ZN(n20582) );
INV_X1 U22517 ( .A(n23395), .ZN(n20504) );
INV_X1 U22518 ( .A(n23402), .ZN(n20542) );
INV_X1 U22519 ( .A(n23411), .ZN(n20580) );
INV_X1 U22520 ( .A(n23545), .ZN(n20502) );
INV_X1 U22521 ( .A(n23552), .ZN(n20540) );
INV_X1 U22522 ( .A(n23561), .ZN(n20578) );
INV_X1 U22523 ( .A(n23707), .ZN(n20538) );
INV_X1 U22524 ( .A(n23716), .ZN(n20576) );
INV_X1 U22525 ( .A(n23871), .ZN(n20536) );
INV_X1 U22526 ( .A(n23880), .ZN(n20574) );
NAND2_X1 U22527 ( .A1(n3745), .A2(n3746), .ZN(n3437) );
NOR2_X1 U22528 ( .A1(n3752), .A2(n3753), .ZN(n3745) );
NOR2_X1 U22529 ( .A1(n3747), .A2(n3748), .ZN(n3746) );
NOR2_X1 U22530 ( .A1(n11507), .A2(n20931), .ZN(n3753) );
NAND2_X1 U22531 ( .A1(n3732), .A2(n3733), .ZN(n3432) );
NOR2_X1 U22532 ( .A1(n3741), .A2(n3742), .ZN(n3732) );
NOR2_X1 U22533 ( .A1(n3734), .A2(n3735), .ZN(n3733) );
NOR2_X1 U22534 ( .A1(n11511), .A2(n20931), .ZN(n3742) );
INV_X1 U22535 ( .A(n23057), .ZN(n20551) );
INV_X1 U22536 ( .A(n23065), .ZN(n20475) );
INV_X1 U22537 ( .A(n23073), .ZN(n20400) );
INV_X1 U22538 ( .A(n23081), .ZN(n20324) );
INV_X1 U22539 ( .A(n22785), .ZN(n20629) );
INV_X1 U22540 ( .A(n22953), .ZN(n20625) );
INV_X1 U22541 ( .A(n22583), .ZN(n20637) );
INV_X1 U22542 ( .A(n22617), .ZN(n20635) );
INV_X1 U22543 ( .A(n22662), .ZN(n20633) );
INV_X1 U22544 ( .A(n22718), .ZN(n20631) );
INV_X1 U22545 ( .A(n22863), .ZN(n20627) );
INV_X1 U22546 ( .A(n23153), .ZN(n20621) );
INV_X1 U22547 ( .A(n23280), .ZN(n20619) );
INV_X1 U22548 ( .A(n23419), .ZN(n20617) );
INV_X1 U22549 ( .A(n23569), .ZN(n20615) );
INV_X1 U22550 ( .A(n23724), .ZN(n20613) );
INV_X1 U22551 ( .A(n23037), .ZN(n20623) );
INV_X1 U22552 ( .A(n23330), .ZN(n20243) );
INV_X1 U22553 ( .A(n23043), .ZN(n20622) );
INV_X1 U22554 ( .A(n23137), .ZN(n20587) );
INV_X1 U22555 ( .A(n23105), .ZN(n20435) );
INV_X1 U22556 ( .A(n23216), .ZN(n20355) );
INV_X1 U22557 ( .A(n23473), .ZN(n20205) );
INV_X1 U22558 ( .A(n22769), .ZN(n20595) );
INV_X1 U22559 ( .A(n22937), .ZN(n20591) );
INV_X1 U22560 ( .A(n23371), .ZN(n20427) );
INV_X1 U22561 ( .A(n23505), .ZN(n20351) );
INV_X1 U22562 ( .A(n23644), .ZN(n20275) );
INV_X1 U22563 ( .A(n24196), .ZN(n20569) );
INV_X1 U22564 ( .A(n22921), .ZN(n20515) );
INV_X1 U22565 ( .A(n23121), .ZN(n20511) );
INV_X1 U22566 ( .A(n23232), .ZN(n20429) );
INV_X1 U22567 ( .A(n23339), .ZN(n20279) );
INV_X1 U22568 ( .A(n23355), .ZN(n20353) );
INV_X1 U22569 ( .A(n23489), .ZN(n20277) );
INV_X1 U22570 ( .A(n23628), .ZN(n20203) );
INV_X1 U22571 ( .A(n23792), .ZN(n20201) );
INV_X1 U22572 ( .A(n22646), .ZN(n20599) );
INV_X1 U22573 ( .A(n22615), .ZN(n20601) );
INV_X1 U22574 ( .A(n22753), .ZN(n20519) );
INV_X1 U22575 ( .A(n22700), .ZN(n20521) );
INV_X1 U22576 ( .A(n22716), .ZN(n20597) );
INV_X1 U22577 ( .A(n22905), .ZN(n20439) );
INV_X1 U22578 ( .A(n22829), .ZN(n20441) );
INV_X1 U22579 ( .A(n22845), .ZN(n20517) );
INV_X1 U22580 ( .A(n22861), .ZN(n20593) );
INV_X1 U22581 ( .A(n23089), .ZN(n20361) );
INV_X1 U22582 ( .A(n23248), .ZN(n20505) );
INV_X1 U22583 ( .A(n23264), .ZN(n20581) );
INV_X1 U22584 ( .A(n23387), .ZN(n20503) );
INV_X1 U22585 ( .A(n23403), .ZN(n20579) );
INV_X1 U22586 ( .A(n23521), .ZN(n20425) );
INV_X1 U22587 ( .A(n23537), .ZN(n20501) );
INV_X1 U22588 ( .A(n23660), .ZN(n20349) );
INV_X1 U22589 ( .A(n23676), .ZN(n20423) );
INV_X1 U22590 ( .A(n23808), .ZN(n20273) );
INV_X1 U22591 ( .A(n23824), .ZN(n20347) );
INV_X1 U22592 ( .A(n23957), .ZN(n20199) );
INV_X1 U22593 ( .A(n23973), .ZN(n20271) );
INV_X1 U22594 ( .A(n24116), .ZN(n20197) );
INV_X1 U22595 ( .A(n24383), .ZN(n20159) );
INV_X1 U22596 ( .A(n23553), .ZN(n20577) );
INV_X1 U22597 ( .A(n23692), .ZN(n20499) );
INV_X1 U22598 ( .A(n23708), .ZN(n20575) );
INV_X1 U22599 ( .A(n23840), .ZN(n20421) );
INV_X1 U22600 ( .A(n23856), .ZN(n20497) );
INV_X1 U22601 ( .A(n23872), .ZN(n20573) );
INV_X1 U22602 ( .A(n23989), .ZN(n20345) );
INV_X1 U22603 ( .A(n24005), .ZN(n20419) );
INV_X1 U22604 ( .A(n24021), .ZN(n20495) );
INV_X1 U22605 ( .A(n24037), .ZN(n20571) );
INV_X1 U22606 ( .A(n24132), .ZN(n20269) );
INV_X1 U22607 ( .A(n24148), .ZN(n20343) );
INV_X1 U22608 ( .A(n24164), .ZN(n20417) );
INV_X1 U22609 ( .A(n24180), .ZN(n20493) );
INV_X1 U22610 ( .A(n24271), .ZN(n20231) );
INV_X1 U22611 ( .A(n24287), .ZN(n20304) );
INV_X1 U22612 ( .A(n24303), .ZN(n20378) );
INV_X1 U22613 ( .A(n24319), .ZN(n20453) );
INV_X1 U22614 ( .A(n24400), .ZN(n20193) );
INV_X1 U22615 ( .A(n24416), .ZN(n20265) );
INV_X1 U22616 ( .A(n24432), .ZN(n20339) );
INV_X1 U22617 ( .A(n24448), .ZN(n20413) );
INV_X1 U22618 ( .A(n24539), .ZN(n20227) );
INV_X1 U22619 ( .A(n24555), .ZN(n20300) );
INV_X1 U22620 ( .A(n24629), .ZN(n20155) );
INV_X1 U22621 ( .A(n24646), .ZN(n20189) );
INV_X1 U22622 ( .A(n22566), .ZN(n20636) );
INV_X1 U22623 ( .A(n22653), .ZN(n20632) );
INV_X1 U22624 ( .A(n22606), .ZN(n20561) );
INV_X1 U22625 ( .A(n22623), .ZN(n20634) );
INV_X1 U22626 ( .A(n22760), .ZN(n20557) );
INV_X1 U22627 ( .A(n22691), .ZN(n20481) );
INV_X1 U22628 ( .A(n22707), .ZN(n20559) );
INV_X1 U22629 ( .A(n22724), .ZN(n20630) );
INV_X1 U22630 ( .A(n22912), .ZN(n20477) );
INV_X1 U22631 ( .A(n22820), .ZN(n20402) );
INV_X1 U22632 ( .A(n22836), .ZN(n20479) );
INV_X1 U22633 ( .A(n22852), .ZN(n20555) );
INV_X1 U22634 ( .A(n22869), .ZN(n20626) );
INV_X1 U22635 ( .A(n23096), .ZN(n20398) );
INV_X1 U22636 ( .A(n23201), .ZN(n20281) );
INV_X1 U22637 ( .A(n23207), .ZN(n20318) );
INV_X1 U22638 ( .A(n23255), .ZN(n20543) );
INV_X1 U22639 ( .A(n23271), .ZN(n20618) );
INV_X1 U22640 ( .A(n23394), .ZN(n20541) );
INV_X1 U22641 ( .A(n23410), .ZN(n20616) );
INV_X1 U22642 ( .A(n23528), .ZN(n20463) );
INV_X1 U22643 ( .A(n23544), .ZN(n20539) );
INV_X1 U22644 ( .A(n23667), .ZN(n20386) );
INV_X1 U22645 ( .A(n23683), .ZN(n20461) );
INV_X1 U22646 ( .A(n23815), .ZN(n20310) );
INV_X1 U22647 ( .A(n23831), .ZN(n20384) );
INV_X1 U22648 ( .A(n23964), .ZN(n20235) );
INV_X1 U22649 ( .A(n23980), .ZN(n20308) );
INV_X1 U22650 ( .A(n24123), .ZN(n20233) );
INV_X1 U22651 ( .A(n24246), .ZN(n20161) );
INV_X1 U22652 ( .A(n23053), .ZN(n20589) );
INV_X1 U22653 ( .A(n23061), .ZN(n20513) );
INV_X1 U22654 ( .A(n23069), .ZN(n20437) );
INV_X1 U22655 ( .A(n23077), .ZN(n20363) );
INV_X1 U22656 ( .A(n23560), .ZN(n20614) );
INV_X1 U22657 ( .A(n23699), .ZN(n20537) );
INV_X1 U22658 ( .A(n23715), .ZN(n20612) );
INV_X1 U22659 ( .A(n23847), .ZN(n20459) );
INV_X1 U22660 ( .A(n23863), .ZN(n20535) );
INV_X1 U22661 ( .A(n23996), .ZN(n20382) );
INV_X1 U22662 ( .A(n24012), .ZN(n20457) );
INV_X1 U22663 ( .A(n24028), .ZN(n20533) );
INV_X1 U22664 ( .A(n24139), .ZN(n20306) );
INV_X1 U22665 ( .A(n24155), .ZN(n20380) );
INV_X1 U22666 ( .A(n24171), .ZN(n20455) );
INV_X1 U22667 ( .A(n24187), .ZN(n20531) );
INV_X1 U22668 ( .A(n24262), .ZN(n20195) );
INV_X1 U22669 ( .A(n24278), .ZN(n20267) );
INV_X1 U22670 ( .A(n24294), .ZN(n20341) );
INV_X1 U22671 ( .A(n24310), .ZN(n20415) );
INV_X1 U22672 ( .A(n24326), .ZN(n20491) );
INV_X1 U22673 ( .A(n24407), .ZN(n20229) );
INV_X1 U22674 ( .A(n24423), .ZN(n20302) );
INV_X1 U22675 ( .A(n24439), .ZN(n20376) );
INV_X1 U22676 ( .A(n24508), .ZN(n20157) );
INV_X1 U22677 ( .A(n24530), .ZN(n20191) );
INV_X1 U22678 ( .A(n24546), .ZN(n20263) );
INV_X1 U22679 ( .A(n24653), .ZN(n20225) );
INV_X1 U22680 ( .A(n24732), .ZN(n20153) );
INV_X1 U22681 ( .A(n22582), .ZN(n20667) );
INV_X1 U22682 ( .A(n22573), .ZN(n20668) );
INV_X1 U22683 ( .A(n22661), .ZN(n20663) );
INV_X1 U22684 ( .A(n22630), .ZN(n20664) );
INV_X1 U22685 ( .A(n22784), .ZN(n20659) );
INV_X1 U22686 ( .A(n22731), .ZN(n20660) );
INV_X1 U22687 ( .A(n22952), .ZN(n20656) );
INV_X1 U22688 ( .A(n22877), .ZN(n20657) );
INV_X1 U22689 ( .A(n23152), .ZN(n20655) );
INV_X1 U22690 ( .A(n23279), .ZN(n20653) );
INV_X1 U22691 ( .A(n23045), .ZN(n20671) );
INV_X1 U22692 ( .A(n23418), .ZN(n20651) );
INV_X1 U22693 ( .A(n23568), .ZN(n20649) );
INV_X1 U22694 ( .A(n24044), .ZN(n20609) );
INV_X1 U22695 ( .A(n23723), .ZN(n20647) );
INV_X1 U22696 ( .A(n23879), .ZN(n20611) );
NAND2_X1 U22697 ( .A1(n5932), .A2(n5933), .ZN(ex_block_i_alu_i_adder_in_b_2) );
NOR2_X1 U22698 ( .A1(n5934), .A2(n5935), .ZN(n5933) );
NOR2_X1 U22699 ( .A1(n5938), .A2(n5939), .ZN(n5932) );
NOR2_X1 U22700 ( .A1(rf_rdata_b_ecc_i_1_), .A2(n20959), .ZN(n5934) );
NAND2_X1 U22701 ( .A1(n5878), .A2(n5879), .ZN(ex_block_i_alu_i_adder_in_b_3) );
NOR2_X1 U22702 ( .A1(n5880), .A2(n5881), .ZN(n5879) );
NOR2_X1 U22703 ( .A1(n5884), .A2(n5885), .ZN(n5878) );
NOR2_X1 U22704 ( .A1(rf_rdata_b_ecc_i_2_), .A2(n20959), .ZN(n5880) );
NAND2_X1 U22705 ( .A1(n5858), .A2(n5859), .ZN(ex_block_i_alu_i_adder_in_b_5) );
NOR2_X1 U22706 ( .A1(n5860), .A2(n5861), .ZN(n5859) );
NOR2_X1 U22707 ( .A1(n5864), .A2(n5865), .ZN(n5858) );
NOR2_X1 U22708 ( .A1(rf_rdata_b_ecc_i_4_), .A2(n20959), .ZN(n5860) );
INV_X1 U22709 ( .A(n25184), .ZN(n20548) );
INV_X1 U22710 ( .A(n22547), .ZN(n20640) );
NAND2_X1 U22711 ( .A1(n10473), .A2(n10474), .ZN(alu_operand_b_ex_4) );
NOR2_X1 U22712 ( .A1(n10475), .A2(n10476), .ZN(n10473) );
NAND2_X1 U22713 ( .A1(rf_rdata_b_ecc_i_4_), .A2(n20950), .ZN(n10474) );
NOR2_X1 U22714 ( .A1(n11311), .A2(n10158), .ZN(n10475) );
INV_X1 U22715 ( .A(n23046), .ZN(n20674) );
INV_X1 U22716 ( .A(n23200), .ZN(n20285) );
INV_X1 U22717 ( .A(n25195), .ZN(n20547) );
INV_X1 U22718 ( .A(n25202), .ZN(n20509) );
INV_X1 U22719 ( .A(n25209), .ZN(n20471) );
INV_X1 U22720 ( .A(n25216), .ZN(n20433) );
INV_X1 U22721 ( .A(n25223), .ZN(n20396) );
INV_X1 U22722 ( .A(n25230), .ZN(n20359) );
INV_X1 U22723 ( .A(n25237), .ZN(n20322) );
INV_X1 U22724 ( .A(n25185), .ZN(n20583) );
INV_X1 U22725 ( .A(n22557), .ZN(n20669) );
INV_X1 U22726 ( .A(n22616), .ZN(n20665) );
INV_X1 U22727 ( .A(n22591), .ZN(n20666) );
INV_X1 U22728 ( .A(n22717), .ZN(n20661) );
INV_X1 U22729 ( .A(n22862), .ZN(n20658) );
INV_X1 U22730 ( .A(n23036), .ZN(n20670) );
INV_X1 U22731 ( .A(n23161), .ZN(n20654) );
INV_X1 U22732 ( .A(n23288), .ZN(n20652) );
INV_X1 U22733 ( .A(n23427), .ZN(n20650) );
INV_X1 U22734 ( .A(n23577), .ZN(n20648) );
NAND2_X1 U22735 ( .A1(n5936), .A2(n5937), .ZN(n5935) );
NAND2_X1 U22736 ( .A1(n20958), .A2(n11164), .ZN(n5937) );
NAND2_X1 U22737 ( .A1(n5818), .A2(n20756), .ZN(n5936) );
NAND2_X1 U22738 ( .A1(n6088), .A2(n6089), .ZN(n6087) );
NAND2_X1 U22739 ( .A1(n20958), .A2(n11165), .ZN(n6089) );
NAND2_X1 U22740 ( .A1(n16410), .A2(n20760), .ZN(n6088) );
NAND2_X1 U22741 ( .A1(n5882), .A2(n5883), .ZN(n5881) );
NAND2_X1 U22742 ( .A1(n20958), .A2(n11163), .ZN(n5883) );
NAND2_X1 U22743 ( .A1(n5818), .A2(n20752), .ZN(n5882) );
NAND2_X1 U22744 ( .A1(n5872), .A2(n5873), .ZN(n5871) );
NAND2_X1 U22745 ( .A1(n20958), .A2(n11162), .ZN(n5873) );
NAND2_X1 U22746 ( .A1(n5818), .A2(n20746), .ZN(n5872) );
NAND2_X1 U22747 ( .A1(n5940), .A2(n5941), .ZN(n5939) );
NAND2_X1 U22748 ( .A1(n11231), .A2(n20960), .ZN(n5941) );
NAND2_X1 U22749 ( .A1(n16409), .A2(n20869), .ZN(n5940) );
NAND2_X1 U22750 ( .A1(n6092), .A2(n6093), .ZN(n6091) );
NAND2_X1 U22751 ( .A1(n11220), .A2(n20960), .ZN(n6093) );
NAND2_X1 U22752 ( .A1(n16409), .A2(n20871), .ZN(n6092) );
NAND2_X1 U22753 ( .A1(n5886), .A2(n5887), .ZN(n5885) );
NAND2_X1 U22754 ( .A1(n11242), .A2(n20960), .ZN(n5887) );
NAND2_X1 U22755 ( .A1(n16409), .A2(n20864), .ZN(n5886) );
NAND2_X1 U22756 ( .A1(n5876), .A2(n5877), .ZN(n5875) );
NAND2_X1 U22757 ( .A1(n11245), .A2(n20960), .ZN(n5877) );
NAND2_X1 U22758 ( .A1(n16409), .A2(n20861), .ZN(n5876) );
INV_X1 U22759 ( .A(n25360), .ZN(n20075) );
INV_X1 U22760 ( .A(n25276), .ZN(n20033) );
INV_X1 U22761 ( .A(n25290), .ZN(n20040) );
INV_X1 U22762 ( .A(n25304), .ZN(n20047) );
INV_X1 U22763 ( .A(n25318), .ZN(n20054) );
INV_X1 U22764 ( .A(n25332), .ZN(n20061) );
INV_X1 U22765 ( .A(n25346), .ZN(n20068) );
INV_X1 U22766 ( .A(n25353), .ZN(n20072) );
INV_X1 U22767 ( .A(n25283), .ZN(n20037) );
INV_X1 U22768 ( .A(n25297), .ZN(n20044) );
INV_X1 U22769 ( .A(n25311), .ZN(n20051) );
INV_X1 U22770 ( .A(n25325), .ZN(n20058) );
INV_X1 U22771 ( .A(n25339), .ZN(n20065) );
INV_X1 U22772 ( .A(n24393), .ZN(n20102) );
INV_X1 U22773 ( .A(n24639), .ZN(n20099) );
AND2_X1 U22774 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_30), .ZN(n434) );
AND2_X1 U22775 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_25), .ZN(n676) );
AND2_X1 U22776 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_26), .ZN(n637) );
AND2_X1 U22777 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_27), .ZN(n597) );
AND2_X1 U22778 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_28), .ZN(n557) );
AND2_X1 U22779 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_29), .ZN(n517) );
INV_X1 U22780 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N63), .ZN(n20039) );
INV_X1 U22781 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N64), .ZN(n20036) );
INV_X1 U22782 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N65), .ZN(n20032) );
INV_X1 U22783 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N66), .ZN(n20027) );
INV_X1 U22784 ( .A(n25245), .ZN(n20073) );
INV_X1 U22785 ( .A(n25247), .ZN(n20066) );
INV_X1 U22786 ( .A(n25243), .ZN(n20083) );
INV_X1 U22787 ( .A(n23953), .ZN(n20082) );
INV_X1 U22788 ( .A(n24112), .ZN(n20077) );
INV_X1 U22789 ( .A(n24396), .ZN(n20070) );
INV_X1 U22790 ( .A(n24642), .ZN(n20063) );
INV_X1 U22791 ( .A(n24113), .ZN(n20076) );
INV_X1 U22792 ( .A(n24397), .ZN(n20069) );
INV_X1 U22793 ( .A(n24643), .ZN(n20062) );
NAND2_X1 U22794 ( .A1(n1751), .A2(n1752), .ZN(instr_addr_o_30_) );
NAND2_X1 U22795 ( .A1(n15929), .A2(n15980), .ZN(n1752) );
NOR2_X1 U22796 ( .A1(n1754), .A2(n1755), .ZN(n1751) );
NOR2_X1 U22797 ( .A1(n10552), .A2(n1706), .ZN(n1755) );
NAND2_X1 U22798 ( .A1(n1745), .A2(n1746), .ZN(instr_addr_o_31_) );
NAND2_X1 U22799 ( .A1(n15929), .A2(n15981), .ZN(n1746) );
NOR2_X1 U22800 ( .A1(n1748), .A2(n1749), .ZN(n1745) );
NOR2_X1 U22801 ( .A1(n10550), .A2(n16459), .ZN(n1749) );
NAND2_X2 U22802 ( .A1(n5623), .A2(n5624), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6) );
NAND2_X1 U22803 ( .A1(rf_rdata_a_ecc_i_6_), .A2(n11299), .ZN(n5623) );
NAND2_X1 U22804 ( .A1(rf_rdata_a_ecc_i_22_), .A2(n5274), .ZN(n5624) );
NAND2_X2 U22805 ( .A1(n5621), .A2(n5622), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7) );
NAND2_X1 U22806 ( .A1(rf_rdata_a_ecc_i_7_), .A2(n11299), .ZN(n5621) );
NAND2_X1 U22807 ( .A1(rf_rdata_a_ecc_i_23_), .A2(n5274), .ZN(n5622) );
NAND2_X2 U22808 ( .A1(n5619), .A2(n5620), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8) );
NAND2_X1 U22809 ( .A1(rf_rdata_a_ecc_i_8_), .A2(n11299), .ZN(n5619) );
NAND2_X1 U22810 ( .A1(rf_rdata_a_ecc_i_24_), .A2(n5274), .ZN(n5620) );
NAND2_X2 U22811 ( .A1(n5617), .A2(n5618), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9) );
NAND2_X1 U22812 ( .A1(n11299), .A2(rf_rdata_a_ecc_i_9_), .ZN(n5617) );
NAND2_X1 U22813 ( .A1(rf_rdata_a_ecc_i_25_), .A2(n5274), .ZN(n5618) );
NAND2_X2 U22814 ( .A1(n5645), .A2(n5646), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10) );
NAND2_X1 U22815 ( .A1(rf_rdata_a_ecc_i_10_), .A2(n11299), .ZN(n5645) );
NAND2_X1 U22816 ( .A1(rf_rdata_a_ecc_i_26_), .A2(n5274), .ZN(n5646) );
NAND2_X1 U22817 ( .A1(n10022), .A2(n15892), .ZN(n10029) );
NAND2_X1 U22818 ( .A1(rf_rdata_b_ecc_i_10_), .A2(n16356), .ZN(n10028) );
NAND2_X1 U22819 ( .A1(n8768), .A2(n8769), .ZN(n240) );
NAND2_X1 U22820 ( .A1(n16366), .A2(crash_dump_o_37_), .ZN(n8769) );
NOR2_X1 U22821 ( .A1(n8771), .A2(n8772), .ZN(n8768) );
NOR2_X1 U22822 ( .A1(n11466), .A2(n8773), .ZN(n8772) );
NAND2_X1 U22823 ( .A1(n9829), .A2(n9830), .ZN(n1295) );
NAND2_X1 U22824 ( .A1(n20947), .A2(crash_dump_o_106_), .ZN(n9830) );
NOR2_X1 U22825 ( .A1(n9831), .A2(n9832), .ZN(n9829) );
NOR2_X1 U22826 ( .A1(n11040), .A2(n8600), .ZN(n9832) );
NAND2_X1 U22827 ( .A1(n8637), .A2(n8638), .ZN(n107) );
NAND2_X1 U22828 ( .A1(n20947), .A2(crash_dump_o_104_), .ZN(n8638) );
NOR2_X1 U22829 ( .A1(n8639), .A2(n8640), .ZN(n8637) );
NOR2_X1 U22830 ( .A1(n11038), .A2(n8600), .ZN(n8640) );
NAND2_X1 U22831 ( .A1(n8595), .A2(n8596), .ZN(n51) );
NAND2_X1 U22832 ( .A1(n20947), .A2(crash_dump_o_105_), .ZN(n8596) );
NOR2_X1 U22833 ( .A1(n8598), .A2(n8599), .ZN(n8595) );
NOR2_X1 U22834 ( .A1(n11039), .A2(n8600), .ZN(n8599) );
NAND2_X1 U22835 ( .A1(n10046), .A2(n10047), .ZN(n149) );
NAND2_X1 U22836 ( .A1(n10022), .A2(n15815), .ZN(n10047) );
NAND2_X1 U22837 ( .A1(rf_rdata_b_ecc_i_7_), .A2(n20950), .ZN(n10046) );
NAND2_X1 U22838 ( .A1(n10023), .A2(n10024), .ZN(n54) );
NAND2_X1 U22839 ( .A1(n10022), .A2(n15918), .ZN(n10024) );
NAND2_X1 U22840 ( .A1(rf_rdata_b_ecc_i_9_), .A2(n20950), .ZN(n10023) ); 
INV_X1 U22841 ( .A(rf_rdata_a_ecc_i_10_), .ZN(n20711) );
INV_X1 U22842 ( .A(rf_rdata_a_ecc_i_9_), .ZN(n20715) );
INV_X1 U22843 ( .A(rf_rdata_a_ecc_i_8_), .ZN(n20719) );
INV_X1 U22844 ( .A(rf_rdata_a_ecc_i_7_), .ZN(n20724) );
INV_X1 U22845 ( .A(rf_rdata_a_ecc_i_6_), .ZN(n20730) );
INV_X1 U22846 ( .A(rf_rdata_a_ecc_i_5_), .ZN(n20735) );
NAND2_X1 U22847 ( .A1(n8726), .A2(n8727), .ZN(n213) );
NAND2_X1 U22848 ( .A1(n20947), .A2(crash_dump_o_102_), .ZN(n8727) );
NOR2_X1 U22849 ( .A1(n8728), .A2(n8729), .ZN(n8726) );
NOR2_X1 U22850 ( .A1(n11036), .A2(n16365), .ZN(n8729) );
NAND2_X1 U22851 ( .A1(n8689), .A2(n8690), .ZN(n170) );
NAND2_X1 U22852 ( .A1(n20947), .A2(crash_dump_o_103_), .ZN(n8690) );
NOR2_X1 U22853 ( .A1(n8691), .A2(n8692), .ZN(n8689) );
NOR2_X1 U22854 ( .A1(n11037), .A2(n16365), .ZN(n8692) );
NAND2_X1 U22855 ( .A1(n5838), .A2(n5839), .ZN(ex_block_i_alu_i_adder_in_b_7) );
NOR2_X1 U22856 ( .A1(n5840), .A2(n5841), .ZN(n5839) );
NOR2_X1 U22857 ( .A1(n5844), .A2(n5845), .ZN(n5838) );
NOR2_X1 U22858 ( .A1(rf_rdata_b_ecc_i_6_), .A2(n20959), .ZN(n5840) );
NAND2_X1 U22859 ( .A1(n5827), .A2(n5828), .ZN(ex_block_i_alu_i_adder_in_b_8) );
NOR2_X1 U22860 ( .A1(n5829), .A2(n5830), .ZN(n5828) );
NOR2_X1 U22861 ( .A1(n5833), .A2(n5834), .ZN(n5827) );
NOR2_X1 U22862 ( .A1(rf_rdata_b_ecc_i_7_), .A2(n20959), .ZN(n5829) );
NAND2_X1 U22863 ( .A1(n6205), .A2(n6206), .ZN(ex_block_i_alu_i_adder_in_b_11) );
NOR2_X1 U22864 ( .A1(n6207), .A2(n6208), .ZN(n6206) );
NOR2_X1 U22865 ( .A1(n6211), .A2(n6212), .ZN(n6205) );
NOR2_X1 U22866 ( .A1(rf_rdata_b_ecc_i_10_), .A2(n20959), .ZN(n6207) );
INV_X1 U22867 ( .A(n22821), .ZN(n20364) );
INV_X1 U22868 ( .A(n22828), .ZN(n20401) );
INV_X1 U22869 ( .A(n22837), .ZN(n20438) );
INV_X1 U22870 ( .A(n22844), .ZN(n20476) );
INV_X1 U22871 ( .A(n22853), .ZN(n20514) );
INV_X1 U22872 ( .A(n24195), .ZN(n20532) );
INV_X1 U22873 ( .A(n24334), .ZN(n20492) );
INV_X1 U22874 ( .A(n24463), .ZN(n20452) );
INV_X1 U22875 ( .A(n22607), .ZN(n20522) );
INV_X1 U22876 ( .A(n22752), .ZN(n20482) );
INV_X1 U22877 ( .A(n22761), .ZN(n20520) );
INV_X1 U22878 ( .A(n22692), .ZN(n20442) );
INV_X1 U22879 ( .A(n22699), .ZN(n20480) );
INV_X1 U22880 ( .A(n22708), .ZN(n20518) );
INV_X1 U22881 ( .A(n22904), .ZN(n20403) );
INV_X1 U22882 ( .A(n22913), .ZN(n20440) );
INV_X1 U22883 ( .A(n22920), .ZN(n20478) );
INV_X1 U22884 ( .A(n23097), .ZN(n20362) );
INV_X1 U22885 ( .A(n23104), .ZN(n20399) );
INV_X1 U22886 ( .A(n23113), .ZN(n20436) );
INV_X1 U22887 ( .A(n23120), .ZN(n20474) );
INV_X1 U22888 ( .A(n23224), .ZN(n20356) );
INV_X1 U22889 ( .A(n23231), .ZN(n20393) );
INV_X1 U22890 ( .A(n23240), .ZN(n20430) );
INV_X1 U22891 ( .A(n23247), .ZN(n20468) );
INV_X1 U22892 ( .A(n23354), .ZN(n20317) );
INV_X1 U22893 ( .A(n23363), .ZN(n20354) );
INV_X1 U22894 ( .A(n23370), .ZN(n20391) );
INV_X1 U22895 ( .A(n23379), .ZN(n20428) );
INV_X1 U22896 ( .A(n23386), .ZN(n20466) );
INV_X1 U22897 ( .A(n23504), .ZN(n20315) );
INV_X1 U22898 ( .A(n23513), .ZN(n20352) );
INV_X1 U22899 ( .A(n23520), .ZN(n20389) );
INV_X1 U22900 ( .A(n23529), .ZN(n20426) );
INV_X1 U22901 ( .A(n23536), .ZN(n20464) );
INV_X1 U22902 ( .A(n23668), .ZN(n20350) );
INV_X1 U22903 ( .A(n23675), .ZN(n20387) );
INV_X1 U22904 ( .A(n23684), .ZN(n20424) );
INV_X1 U22905 ( .A(n23691), .ZN(n20462) );
INV_X1 U22906 ( .A(n23700), .ZN(n20500) );
INV_X1 U22907 ( .A(n23832), .ZN(n20348) );
INV_X1 U22908 ( .A(n23839), .ZN(n20385) );
INV_X1 U22909 ( .A(n23848), .ZN(n20422) );
INV_X1 U22910 ( .A(n23855), .ZN(n20460) );
INV_X1 U22911 ( .A(n23864), .ZN(n20498) );
INV_X1 U22912 ( .A(n24004), .ZN(n20383) );
INV_X1 U22913 ( .A(n24013), .ZN(n20420) );
INV_X1 U22914 ( .A(n24020), .ZN(n20458) );
INV_X1 U22915 ( .A(n24029), .ZN(n20496) );
INV_X1 U22916 ( .A(n24036), .ZN(n20534) );
INV_X1 U22917 ( .A(n24163), .ZN(n20381) );
INV_X1 U22918 ( .A(n24172), .ZN(n20418) );
INV_X1 U22919 ( .A(n24179), .ZN(n20456) );
INV_X1 U22920 ( .A(n24188), .ZN(n20494) );
INV_X1 U22921 ( .A(n24318), .ZN(n20416) );
INV_X1 U22922 ( .A(n24327), .ZN(n20454) );
NAND2_X1 U22923 ( .A1(n3818), .A2(n3819), .ZN(n3472) );
NOR2_X1 U22924 ( .A1(n3825), .A2(n3826), .ZN(n3818) );
NOR2_X1 U22925 ( .A1(n3820), .A2(n3821), .ZN(n3819) );
NOR2_X1 U22926 ( .A1(n10932), .A2(n20931), .ZN(n3826) );
NAND2_X1 U22927 ( .A1(n3795), .A2(n3796), .ZN(n3462) );
NOR2_X1 U22928 ( .A1(n3802), .A2(n3803), .ZN(n3795) );
NOR2_X1 U22929 ( .A1(n3797), .A2(n3798), .ZN(n3796) );
NOR2_X1 U22930 ( .A1(n10962), .A2(n16355), .ZN(n3803) );
NAND2_X1 U22931 ( .A1(n3756), .A2(n3757), .ZN(n3447) );
NOR2_X1 U22932 ( .A1(n3763), .A2(n3764), .ZN(n3756) );
NOR2_X1 U22933 ( .A1(n3758), .A2(n3759), .ZN(n3757) );
NOR2_X1 U22934 ( .A1(n10624), .A2(n20931), .ZN(n3764) );
INV_X1 U22935 ( .A(n24205), .ZN(n20570) );
INV_X1 U22936 ( .A(n24344), .ZN(n20530) );
INV_X1 U22937 ( .A(n24335), .ZN(n20529) );
INV_X1 U22938 ( .A(n24464), .ZN(n20489) );
INV_X1 U22939 ( .A(n24587), .ZN(n20449) );
INV_X1 U22940 ( .A(n24694), .ZN(n20409) );
INV_X1 U22941 ( .A(n24571), .ZN(n20374) );
INV_X1 U22942 ( .A(n24662), .ZN(n20261) );
INV_X1 U22943 ( .A(n24678), .ZN(n20335) );
INV_X1 U22944 ( .A(n24757), .ZN(n20223) );
INV_X1 U22945 ( .A(n24773), .ZN(n20296) );
INV_X1 U22946 ( .A(n24825), .ZN(n20151) );
INV_X1 U22947 ( .A(n24842), .ZN(n20185) );
INV_X1 U22948 ( .A(n24858), .ZN(n20257) );
INV_X1 U22949 ( .A(n24977), .ZN(n20147) );
INV_X1 U22950 ( .A(n24054), .ZN(n20610) );
INV_X1 U22951 ( .A(n24455), .ZN(n20451) );
INV_X1 U22952 ( .A(n24562), .ZN(n20337) );
INV_X1 U22953 ( .A(n24578), .ZN(n20411) );
INV_X1 U22954 ( .A(n24669), .ZN(n20298) );
INV_X1 U22955 ( .A(n24685), .ZN(n20372) );
INV_X1 U22956 ( .A(n24748), .ZN(n20187) );
INV_X1 U22957 ( .A(n24764), .ZN(n20259) );
INV_X1 U22958 ( .A(n24780), .ZN(n20333) );
INV_X1 U22959 ( .A(n24849), .ZN(n20221) );
INV_X1 U22960 ( .A(n24865), .ZN(n20294) );
INV_X1 U22961 ( .A(n24906), .ZN(n20149) );
INV_X1 U22962 ( .A(n24922), .ZN(n20183) );
NAND2_X1 U22963 ( .A1(n5848), .A2(n5849), .ZN(ex_block_i_alu_i_adder_in_b_6) );
NOR2_X1 U22964 ( .A1(n5850), .A2(n5851), .ZN(n5849) );
NOR2_X1 U22965 ( .A1(n5854), .A2(n5855), .ZN(n5848) );
NOR2_X1 U22966 ( .A1(rf_rdata_b_ecc_i_5_), .A2(n20959), .ZN(n5850) );
NAND2_X1 U22967 ( .A1(n5811), .A2(n5812), .ZN(ex_block_i_alu_i_adder_in_b_9) );
NOR2_X1 U22968 ( .A1(n5813), .A2(n5814), .ZN(n5812) );
NOR2_X1 U22969 ( .A1(n5820), .A2(n5821), .ZN(n5811) );
NOR2_X1 U22970 ( .A1(rf_rdata_b_ecc_i_8_), .A2(n20959), .ZN(n5813) );
NAND2_X1 U22971 ( .A1(n6216), .A2(n6217), .ZN(ex_block_i_alu_i_adder_in_b_10) );
NOR2_X1 U22972 ( .A1(n6218), .A2(n6219), .ZN(n6217) );
NOR2_X1 U22973 ( .A1(n6223), .A2(n6224), .ZN(n6216) );
NOR2_X1 U22974 ( .A1(rf_rdata_b_ecc_i_9_), .A2(n20959), .ZN(n6218) );
INV_X1 U22975 ( .A(n25194), .ZN(n20510) );
INV_X1 U22976 ( .A(n25201), .ZN(n20472) );
INV_X1 U22977 ( .A(n25208), .ZN(n20434) );
INV_X1 U22978 ( .A(n25215), .ZN(n20397) );
NAND2_X1 U22979 ( .A1(n10061), .A2(n10062), .ZN(n255) );
NAND2_X1 U22980 ( .A1(n10022), .A2(n15807), .ZN(n10062) );
NAND2_X1 U22981 ( .A1(rf_rdata_b_ecc_i_5_), .A2(n16356), .ZN(n10061) );
NAND2_X1 U22982 ( .A1(n10020), .A2(n10021), .ZN(n109) );
NAND2_X1 U22983 ( .A1(n10022), .A2(n15982), .ZN(n10021) );
NAND2_X1 U22984 ( .A1(rf_rdata_b_ecc_i_8_), .A2(n20950), .ZN(n10020) );
NAND2_X1 U22985 ( .A1(n10041), .A2(n10042), .ZN(n197) );
NAND2_X1 U22986 ( .A1(n10022), .A2(n15824), .ZN(n10042) );
NAND2_X1 U22987 ( .A1(rf_rdata_b_ecc_i_6_), .A2(n16356), .ZN(n10041) );
NAND2_X1 U22988 ( .A1(n5822), .A2(n5823), .ZN(n5821) );
NAND2_X1 U22989 ( .A1(n11250), .A2(n20960), .ZN(n5823) );
NAND2_X1 U22990 ( .A1(n20835), .A2(n5826), .ZN(n5822) );
NAND2_X1 U22991 ( .A1(n6213), .A2(n6214), .ZN(n6212) );
NAND2_X1 U22992 ( .A1(n11221), .A2(n20960), .ZN(n6214) );
NAND2_X1 U22993 ( .A1(n20830), .A2(n16409), .ZN(n6213) );
NAND2_X1 U22994 ( .A1(n5862), .A2(n5863), .ZN(n5861) );
NAND2_X1 U22995 ( .A1(n20958), .A2(n11161), .ZN(n5863) );
NAND2_X1 U22996 ( .A1(n5818), .A2(n20741), .ZN(n5862) );
NAND2_X1 U22997 ( .A1(n5852), .A2(n5853), .ZN(n5851) );
NAND2_X1 U22998 ( .A1(n20958), .A2(n11160), .ZN(n5853) );
NAND2_X1 U22999 ( .A1(n5818), .A2(n20735), .ZN(n5852) );
NAND2_X1 U23000 ( .A1(n5842), .A2(n5843), .ZN(n5841) );
NAND2_X1 U23001 ( .A1(n20958), .A2(n11159), .ZN(n5843) );
NAND2_X1 U23002 ( .A1(n5818), .A2(n20730), .ZN(n5842) );
NAND2_X1 U23003 ( .A1(n5831), .A2(n5832), .ZN(n5830) );
NAND2_X1 U23004 ( .A1(n20958), .A2(n11158), .ZN(n5832) );
NAND2_X1 U23005 ( .A1(n5818), .A2(n20724), .ZN(n5831) );
NAND2_X1 U23006 ( .A1(n5815), .A2(n5816), .ZN(n5814) );
NAND2_X1 U23007 ( .A1(n20958), .A2(n11157), .ZN(n5816) );
NAND2_X1 U23008 ( .A1(n5818), .A2(n20719), .ZN(n5815) );
NAND2_X1 U23009 ( .A1(n6220), .A2(n6221), .ZN(n6219) );
NAND2_X1 U23010 ( .A1(n20958), .A2(n11156), .ZN(n6221) );
NAND2_X1 U23011 ( .A1(n16410), .A2(n20715), .ZN(n6220) );
NAND2_X1 U23012 ( .A1(n5856), .A2(n5857), .ZN(n5855) );
NAND2_X1 U23013 ( .A1(n11247), .A2(n20960), .ZN(n5857) );
NAND2_X1 U23014 ( .A1(n20846), .A2(n16409), .ZN(n5856) );
NAND2_X1 U23015 ( .A1(n5846), .A2(n5847), .ZN(n5845) );
NAND2_X1 U23016 ( .A1(n11248), .A2(n20960), .ZN(n5847) );
NAND2_X1 U23017 ( .A1(n20841), .A2(n5826), .ZN(n5846) );
NAND2_X1 U23018 ( .A1(n5835), .A2(n5836), .ZN(n5834) );
NAND2_X1 U23019 ( .A1(n11249), .A2(n20960), .ZN(n5836) );
NAND2_X1 U23020 ( .A1(n20839), .A2(n16409), .ZN(n5835) );
NAND2_X1 U23021 ( .A1(n6225), .A2(n6226), .ZN(n6224) );
NAND2_X1 U23022 ( .A1(n11251), .A2(n20960), .ZN(n6226) );
NAND2_X1 U23023 ( .A1(n20833), .A2(n5826), .ZN(n6225) );
INV_X1 U23024 ( .A(n24835), .ZN(n20096) );
INV_X1 U23025 ( .A(n24987), .ZN(n20093) );
AND2_X1 U23026 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_19), .ZN(n947) );
AND2_X1 U23027 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_20), .ZN(n866) );
AND2_X1 U23028 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_21), .ZN(n827) );
AND2_X1 U23029 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_22), .ZN(n789) );
AND2_X1 U23030 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_23), .ZN(n751) );
AND2_X1 U23031 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_24), .ZN(n714) );
INV_X1 U23032 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N54), .ZN(n20071) );
INV_X1 U23033 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N55), .ZN(n20067) );
INV_X1 U23034 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N56), .ZN(n20064) );
INV_X1 U23035 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N57), .ZN(n20060) );
INV_X1 U23036 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N58), .ZN(n20057) );
INV_X1 U23037 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N59), .ZN(n20053) );
INV_X1 U23038 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N60), .ZN(n20050) );
INV_X1 U23039 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N61), .ZN(n20046) );
INV_X1 U23040 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N62), .ZN(n20043) );
INV_X1 U23041 ( .A(n25249), .ZN(n20059) );
INV_X1 U23042 ( .A(n25251), .ZN(n20052) );
INV_X1 U23043 ( .A(n24838), .ZN(n20056) );
INV_X1 U23044 ( .A(n24990), .ZN(n20049) );
INV_X1 U23045 ( .A(n24839), .ZN(n20055) );
INV_X1 U23046 ( .A(n24991), .ZN(n20048) );
NAND2_X1 U23047 ( .A1(n1793), .A2(n1794), .ZN(instr_addr_o_24_) );
NAND2_X1 U23048 ( .A1(n15929), .A2(n15983), .ZN(n1794) );
NOR2_X1 U23049 ( .A1(n1796), .A2(n1797), .ZN(n1793) );
NOR2_X1 U23050 ( .A1(n10564), .A2(n1706), .ZN(n1797) );
NAND2_X1 U23051 ( .A1(n1787), .A2(n1788), .ZN(instr_addr_o_25_) );
NAND2_X1 U23052 ( .A1(n15929), .A2(n16054), .ZN(n1788) );
NOR2_X1 U23053 ( .A1(n1790), .A2(n1791), .ZN(n1787) );
NOR2_X1 U23054 ( .A1(n10562), .A2(n1706), .ZN(n1791) );
NAND2_X1 U23055 ( .A1(n1781), .A2(n1782), .ZN(instr_addr_o_26_) );
NAND2_X1 U23056 ( .A1(n15929), .A2(n15984), .ZN(n1782) );
NOR2_X1 U23057 ( .A1(n1784), .A2(n1785), .ZN(n1781) );
NOR2_X1 U23058 ( .A1(n10560), .A2(n1706), .ZN(n1785) );
NAND2_X1 U23059 ( .A1(n1775), .A2(n1776), .ZN(instr_addr_o_27_) );
NAND2_X1 U23060 ( .A1(n15929), .A2(n16055), .ZN(n1776) );
NOR2_X1 U23061 ( .A1(n1778), .A2(n1779), .ZN(n1775) );
NOR2_X1 U23062 ( .A1(n10558), .A2(n1706), .ZN(n1779) );
NAND2_X1 U23063 ( .A1(n1769), .A2(n1770), .ZN(instr_addr_o_28_) );
NAND2_X1 U23064 ( .A1(n15929), .A2(n16056), .ZN(n1770) );
NOR2_X1 U23065 ( .A1(n1772), .A2(n1773), .ZN(n1769) );
NOR2_X1 U23066 ( .A1(n10556), .A2(n16459), .ZN(n1773) );
NAND2_X1 U23067 ( .A1(n1763), .A2(n1764), .ZN(instr_addr_o_29_) );
NAND2_X1 U23068 ( .A1(n15929), .A2(n15985), .ZN(n1764) );
NOR2_X1 U23069 ( .A1(n1766), .A2(n1767), .ZN(n1763) );
NOR2_X1 U23070 ( .A1(n10554), .A2(n16459), .ZN(n1767) );
NAND2_X2 U23071 ( .A1(n5643), .A2(n5644), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11) );
NAND2_X1 U23072 ( .A1(rf_rdata_a_ecc_i_11_), .A2(n11299), .ZN(n5643) );
NAND2_X1 U23073 ( .A1(rf_rdata_a_ecc_i_27_), .A2(n5274), .ZN(n5644) );
NAND2_X2 U23074 ( .A1(n5641), .A2(n5642), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12) );
NAND2_X1 U23075 ( .A1(rf_rdata_a_ecc_i_12_), .A2(n11299), .ZN(n5641) );
NAND2_X1 U23076 ( .A1(rf_rdata_a_ecc_i_28_), .A2(n5274), .ZN(n5642) );
NAND2_X2 U23077 ( .A1(n5639), .A2(n5640), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13) );
NAND2_X1 U23078 ( .A1(rf_rdata_a_ecc_i_13_), .A2(n11299), .ZN(n5639) );
NAND2_X1 U23079 ( .A1(rf_rdata_a_ecc_i_29_), .A2(n5274), .ZN(n5640) );
NAND2_X2 U23080 ( .A1(n5637), .A2(n5638), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14) );
NAND2_X1 U23081 ( .A1(rf_rdata_a_ecc_i_14_), .A2(n11299), .ZN(n5637) );
NAND2_X1 U23082 ( .A1(rf_rdata_a_ecc_i_30_), .A2(n5274), .ZN(n5638) );
NAND2_X1 U23083 ( .A1(n9592), .A2(n9593), .ZN(n1046) );
NAND2_X1 U23084 ( .A1(n20947), .A2(crash_dump_o_112_), .ZN(n9593) );
NOR2_X1 U23085 ( .A1(n9594), .A2(n9595), .ZN(n9592) );
NOR2_X1 U23086 ( .A1(n11046), .A2(n8600), .ZN(n9595) );
NAND2_X1 U23087 ( .A1(n9630), .A2(n9631), .ZN(n1102) );
NAND2_X1 U23088 ( .A1(n20947), .A2(crash_dump_o_111_), .ZN(n9631) );
NOR2_X1 U23089 ( .A1(n9632), .A2(n9633), .ZN(n9630) );
NOR2_X1 U23090 ( .A1(n11045), .A2(n16365), .ZN(n9633) );
NAND2_X1 U23091 ( .A1(n9792), .A2(n9793), .ZN(n1258) );
NAND2_X1 U23092 ( .A1(n16366), .A2(crash_dump_o_43_), .ZN(n9793) );
NOR2_X1 U23093 ( .A1(n9794), .A2(n9795), .ZN(n9792) );
NOR2_X1 U23094 ( .A1(n11307), .A2(n8773), .ZN(n9795) );
NAND2_X1 U23095 ( .A1(n9667), .A2(n9668), .ZN(n1139) );
NAND2_X1 U23096 ( .A1(n20947), .A2(crash_dump_o_110_), .ZN(n9668) );
NOR2_X1 U23097 ( .A1(n9669), .A2(n9670), .ZN(n9667) );
NOR2_X1 U23098 ( .A1(n11044), .A2(n8600), .ZN(n9670) );
NAND2_X1 U23099 ( .A1(n9704), .A2(n9705), .ZN(n1178) );
NAND2_X1 U23100 ( .A1(n20947), .A2(crash_dump_o_109_), .ZN(n9705) );
NOR2_X1 U23101 ( .A1(n9706), .A2(n9707), .ZN(n9704) );
NOR2_X1 U23102 ( .A1(n11043), .A2(n16365), .ZN(n9707) );
NAND2_X1 U23103 ( .A1(n9744), .A2(n9745), .ZN(n1217) );
NAND2_X1 U23104 ( .A1(n20947), .A2(crash_dump_o_108_), .ZN(n9745) );
NOR2_X1 U23105 ( .A1(n9746), .A2(n9747), .ZN(n9744) );
NOR2_X1 U23106 ( .A1(n11042), .A2(n8600), .ZN(n9747) );
INV_X1 U23107 ( .A(rf_rdata_b_ecc_i_15_), .ZN(n20811) );
INV_X1 U23108 ( .A(rf_rdata_b_ecc_i_14_), .ZN(n20813) );
INV_X1 U23109 ( .A(rf_rdata_b_ecc_i_13_), .ZN(n20815) );
INV_X1 U23110 ( .A(rf_rdata_b_ecc_i_12_), .ZN(n20817) );
NAND2_X1 U23111 ( .A1(n6183), .A2(n6184), .ZN(n1219) );
NOR2_X1 U23112 ( .A1(n6077), .A2(n6185), .ZN(n6183) );
NAND2_X1 U23113 ( .A1(rf_rdata_b_ecc_i_12_), .A2(n20950), .ZN(n6184) );
NOR2_X1 U23114 ( .A1(n11313), .A2(n6079), .ZN(n6185) );
NAND2_X1 U23115 ( .A1(n6169), .A2(n6170), .ZN(n1180) );
NOR2_X1 U23116 ( .A1(n6077), .A2(n6171), .ZN(n6169) );
NAND2_X1 U23117 ( .A1(rf_rdata_b_ecc_i_13_), .A2(n20950), .ZN(n6170) );
NOR2_X1 U23118 ( .A1(n11320), .A2(n6079), .ZN(n6171) );
NAND2_X1 U23119 ( .A1(n6155), .A2(n6156), .ZN(n1141) );
NOR2_X1 U23120 ( .A1(n6077), .A2(n6157), .ZN(n6155) );
NAND2_X1 U23121 ( .A1(rf_rdata_b_ecc_i_14_), .A2(n20950), .ZN(n6156) );
NOR2_X1 U23122 ( .A1(n11329), .A2(n6079), .ZN(n6157) );
INV_X1 U23123 ( .A(rf_rdata_a_ecc_i_11_), .ZN(n20707) );
INV_X1 U23124 ( .A(rf_rdata_a_ecc_i_14_), .ZN(n20695) );
INV_X1 U23125 ( .A(rf_rdata_a_ecc_i_15_), .ZN(n20691) );
INV_X1 U23126 ( .A(rf_rdata_a_ecc_i_16_), .ZN(n20687) );
INV_X1 U23127 ( .A(rf_rdata_a_ecc_i_13_), .ZN(n20699) );
INV_X1 U23128 ( .A(rf_rdata_a_ecc_i_12_), .ZN(n20703) );
NAND2_X1 U23129 ( .A1(n6141), .A2(n6142), .ZN(n1100) );
NOR2_X1 U23130 ( .A1(n6077), .A2(n6143), .ZN(n6141) );
NAND2_X1 U23131 ( .A1(rf_rdata_b_ecc_i_15_), .A2(n20950), .ZN(n6142) );
NOR2_X1 U23132 ( .A1(n6079), .A2(n15890), .ZN(n6143) );
NAND2_X1 U23133 ( .A1(n6128), .A2(n6129), .ZN(n1044) );
NOR2_X1 U23134 ( .A1(n6077), .A2(n6130), .ZN(n6128) );
NAND2_X1 U23135 ( .A1(rf_rdata_b_ecc_i_16_), .A2(n16356), .ZN(n6129) );
NOR2_X1 U23136 ( .A1(n6079), .A2(n15809), .ZN(n6130) );
INV_X1 U23137 ( .A(n23088), .ZN(n20325) );
INV_X1 U23138 ( .A(n23208), .ZN(n20282) );
INV_X1 U23139 ( .A(n23331), .ZN(n20209) );
INV_X1 U23140 ( .A(n23338), .ZN(n20244) );
INV_X1 U23141 ( .A(n23481), .ZN(n20206) );
INV_X1 U23142 ( .A(n23627), .ZN(n20168) );
INV_X1 U23143 ( .A(n24586), .ZN(n20412) );
INV_X1 U23144 ( .A(n24693), .ZN(n20373) );
INV_X1 U23145 ( .A(n23215), .ZN(n20319) );
INV_X1 U23146 ( .A(n23347), .ZN(n20280) );
INV_X1 U23147 ( .A(n23488), .ZN(n20242) );
INV_X1 U23148 ( .A(n23497), .ZN(n20278) );
INV_X1 U23149 ( .A(n23636), .ZN(n20204) );
INV_X1 U23150 ( .A(n23643), .ZN(n20240) );
INV_X1 U23151 ( .A(n23652), .ZN(n20276) );
INV_X1 U23152 ( .A(n23659), .ZN(n20313) );
INV_X1 U23153 ( .A(n23791), .ZN(n20166) );
INV_X1 U23154 ( .A(n23800), .ZN(n20202) );
INV_X1 U23155 ( .A(n23807), .ZN(n20238) );
INV_X1 U23156 ( .A(n23816), .ZN(n20274) );
INV_X1 U23157 ( .A(n23823), .ZN(n20311) );
INV_X1 U23158 ( .A(n23956), .ZN(n20164) );
INV_X1 U23159 ( .A(n23965), .ZN(n20200) );
INV_X1 U23160 ( .A(n23972), .ZN(n20236) );
INV_X1 U23161 ( .A(n23981), .ZN(n20272) );
INV_X1 U23162 ( .A(n23988), .ZN(n20309) );
INV_X1 U23163 ( .A(n23997), .ZN(n20346) );
INV_X1 U23164 ( .A(n24124), .ZN(n20198) );
INV_X1 U23165 ( .A(n24131), .ZN(n20234) );
INV_X1 U23166 ( .A(n24140), .ZN(n20270) );
INV_X1 U23167 ( .A(n24147), .ZN(n20307) );
INV_X1 U23168 ( .A(n24156), .ZN(n20344) );
INV_X1 U23169 ( .A(n24279), .ZN(n20232) );
INV_X1 U23170 ( .A(n24286), .ZN(n20268) );
INV_X1 U23171 ( .A(n24295), .ZN(n20305) );
INV_X1 U23172 ( .A(n24302), .ZN(n20342) );
INV_X1 U23173 ( .A(n24311), .ZN(n20379) );
INV_X1 U23174 ( .A(n24415), .ZN(n20230) );
INV_X1 U23175 ( .A(n24424), .ZN(n20266) );
INV_X1 U23176 ( .A(n24431), .ZN(n20303) );
INV_X1 U23177 ( .A(n24440), .ZN(n20340) );
INV_X1 U23178 ( .A(n24447), .ZN(n20377) );
INV_X1 U23179 ( .A(n24456), .ZN(n20414) );
INV_X1 U23180 ( .A(n24563), .ZN(n20301) );
INV_X1 U23181 ( .A(n24570), .ZN(n20338) );
INV_X1 U23182 ( .A(n24579), .ZN(n20375) );
INV_X1 U23183 ( .A(n24677), .ZN(n20299) );
INV_X1 U23184 ( .A(n24686), .ZN(n20336) );
NAND2_X1 U23185 ( .A1(n3885), .A2(n3886), .ZN(n3513) );
NOR2_X1 U23186 ( .A1(n3892), .A2(n3893), .ZN(n3885) );
NOR2_X1 U23187 ( .A1(n3887), .A2(n3888), .ZN(n3886) );
NOR2_X1 U23188 ( .A1(n10857), .A2(n16355), .ZN(n3893) );
NAND2_X1 U23189 ( .A1(n3874), .A2(n3875), .ZN(n3508) );
NOR2_X1 U23190 ( .A1(n3881), .A2(n3882), .ZN(n3874) );
NOR2_X1 U23191 ( .A1(n3876), .A2(n3877), .ZN(n3875) );
NOR2_X1 U23192 ( .A1(n10872), .A2(n16355), .ZN(n3882) );
NAND2_X1 U23193 ( .A1(n3851), .A2(n3852), .ZN(n3487) );
NOR2_X1 U23194 ( .A1(n3858), .A2(n3859), .ZN(n3851) );
NOR2_X1 U23195 ( .A1(n3853), .A2(n3854), .ZN(n3852) );
NOR2_X1 U23196 ( .A1(n11497), .A2(n20931), .ZN(n3859) );
NAND2_X1 U23197 ( .A1(n3840), .A2(n3841), .ZN(n3482) );
NOR2_X1 U23198 ( .A1(n3847), .A2(n3848), .ZN(n3840) );
NOR2_X1 U23199 ( .A1(n3842), .A2(n3843), .ZN(n3841) );
NOR2_X1 U23200 ( .A1(n10902), .A2(n16355), .ZN(n3848) );
NAND2_X1 U23201 ( .A1(n3829), .A2(n3830), .ZN(n3477) );
NOR2_X1 U23202 ( .A1(n3836), .A2(n3837), .ZN(n3829) );
NOR2_X1 U23203 ( .A1(n3831), .A2(n3832), .ZN(n3830) );
NOR2_X1 U23204 ( .A1(n10917), .A2(n20931), .ZN(n3837) );
INV_X1 U23205 ( .A(n24473), .ZN(n20490) );
INV_X1 U23206 ( .A(n24596), .ZN(n20450) );
INV_X1 U23207 ( .A(n24703), .ZN(n20410) );
INV_X1 U23208 ( .A(n24789), .ZN(n20370) );
INV_X1 U23209 ( .A(n24874), .ZN(n20331) );
INV_X1 U23210 ( .A(n24947), .ZN(n20292) );
INV_X1 U23211 ( .A(n25010), .ZN(n20253) );
INV_X1 U23212 ( .A(n24931), .ZN(n20219) );
INV_X1 U23213 ( .A(n24994), .ZN(n20181) );
INV_X1 U23214 ( .A(n25085), .ZN(n20143) );
INV_X1 U23215 ( .A(n24938), .ZN(n20255) );
INV_X1 U23216 ( .A(n25001), .ZN(n20217) );
INV_X1 U23217 ( .A(n25036), .ZN(n20145) );
INV_X1 U23218 ( .A(n25052), .ZN(n20179) );
INV_X1 U23219 ( .A(n25122), .ZN(n20141) );
NAND2_X1 U23220 ( .A1(n6195), .A2(n6196), .ZN(ex_block_i_alu_i_adder_in_b_12) );
NOR2_X1 U23221 ( .A1(n6197), .A2(n6198), .ZN(n6196) );
NOR2_X1 U23222 ( .A1(n6201), .A2(n6202), .ZN(n6195) );
NOR2_X1 U23223 ( .A1(rf_rdata_b_ecc_i_11_), .A2(n20959), .ZN(n6197) );
INV_X1 U23224 ( .A(n23085), .ZN(n20247) );
INV_X1 U23225 ( .A(n25222), .ZN(n20360) );
INV_X1 U23226 ( .A(n25229), .ZN(n20323) );
INV_X1 U23227 ( .A(n25236), .ZN(n20286) );
NAND2_X1 U23228 ( .A1(n10048), .A2(n10049), .ZN(n1256) );
NAND2_X1 U23229 ( .A1(n10050), .A2(n10051), .ZN(n10049) );
NAND2_X1 U23230 ( .A1(rf_rdata_b_ecc_i_11_), .A2(n20950), .ZN(n10048) );
NAND2_X1 U23231 ( .A1(n10052), .A2(n10053), .ZN(n10050) );
INV_X1 U23232 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_13), .ZN(n20207) );
INV_X1 U23233 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_14), .ZN(n20169) );
NAND2_X1 U23234 ( .A1(n6209), .A2(n6210), .ZN(n6208) );
NAND2_X1 U23235 ( .A1(n20958), .A2(n11218), .ZN(n6210) );
NAND2_X1 U23236 ( .A1(n16410), .A2(n20711), .ZN(n6209) );
NAND2_X1 U23237 ( .A1(n6199), .A2(n6200), .ZN(n6198) );
NAND2_X1 U23238 ( .A1(n20958), .A2(n11186), .ZN(n6200) );
NAND2_X1 U23239 ( .A1(n16410), .A2(n20707), .ZN(n6199) );
NAND2_X1 U23240 ( .A1(n6203), .A2(n6204), .ZN(n6202) );
NAND2_X1 U23241 ( .A1(n11222), .A2(n20960), .ZN(n6204) );
NAND2_X1 U23242 ( .A1(n20828), .A2(n16409), .ZN(n6203) );
INV_X1 U23243 ( .A(n25095), .ZN(n20090) );
AND2_X1 U23244 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_16), .ZN(n1082) );
AND2_X1 U23245 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_17), .ZN(n1024) );
AND2_X1 U23246 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_18), .ZN(n986) );
INV_X1 U23247 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_15), .ZN(n20107) );
INV_X1 U23248 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N49), .ZN(n20170) );
INV_X1 U23249 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N51), .ZN(n20026) );
INV_X1 U23250 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N53), .ZN(n20074) );
INV_X1 U23251 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N52), .ZN(n20078) );
INV_X1 U23252 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N48), .ZN(n20208) );
INV_X1 U23253 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N50), .ZN(n20108) );
INV_X1 U23254 ( .A(n25253), .ZN(n20045) );
INV_X1 U23255 ( .A(n25098), .ZN(n20042) );
INV_X1 U23256 ( .A(n25099), .ZN(n20041) );
NAND2_X1 U23257 ( .A1(n1829), .A2(n1830), .ZN(instr_addr_o_18_) );
NAND2_X1 U23258 ( .A1(n15929), .A2(n15986), .ZN(n1830) );
NOR2_X1 U23259 ( .A1(n1832), .A2(n1833), .ZN(n1829) );
NOR2_X1 U23260 ( .A1(n10576), .A2(n1706), .ZN(n1833) );
NAND2_X1 U23261 ( .A1(n1823), .A2(n1824), .ZN(instr_addr_o_19_) );
NAND2_X1 U23262 ( .A1(n15929), .A2(n15987), .ZN(n1824) );
NOR2_X1 U23263 ( .A1(n1826), .A2(n1827), .ZN(n1823) );
NOR2_X1 U23264 ( .A1(n10574), .A2(n1706), .ZN(n1827) );
NAND2_X1 U23265 ( .A1(n1817), .A2(n1818), .ZN(instr_addr_o_20_) );
NAND2_X1 U23266 ( .A1(n15929), .A2(n16053), .ZN(n1818) );
NOR2_X1 U23267 ( .A1(n1820), .A2(n1821), .ZN(n1817) );
NOR2_X1 U23268 ( .A1(n10572), .A2(n1706), .ZN(n1821) );
NAND2_X1 U23269 ( .A1(n1811), .A2(n1812), .ZN(instr_addr_o_21_) );
NAND2_X1 U23270 ( .A1(n15929), .A2(n15988), .ZN(n1812) );
NOR2_X1 U23271 ( .A1(n1814), .A2(n1815), .ZN(n1811) );
NOR2_X1 U23272 ( .A1(n10570), .A2(n1706), .ZN(n1815) );
NAND2_X1 U23273 ( .A1(n1805), .A2(n1806), .ZN(instr_addr_o_22_) );
NAND2_X1 U23274 ( .A1(n15929), .A2(n15989), .ZN(n1806) );
NOR2_X1 U23275 ( .A1(n1808), .A2(n1809), .ZN(n1805) );
NOR2_X1 U23276 ( .A1(n10568), .A2(n1706), .ZN(n1809) );
NAND2_X1 U23277 ( .A1(n1799), .A2(n1800), .ZN(instr_addr_o_23_) );
NAND2_X1 U23278 ( .A1(n15929), .A2(n15990), .ZN(n1800) );
NOR2_X1 U23279 ( .A1(n1802), .A2(n1803), .ZN(n1799) );
NOR2_X1 U23280 ( .A1(n10566), .A2(n1706), .ZN(n1803) );
NAND2_X2 U23281 ( .A1(n5635), .A2(n5636), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15) );
NAND2_X1 U23282 ( .A1(rf_rdata_a_ecc_i_15_), .A2(n11299), .ZN(n5635) );
NAND2_X1 U23283 ( .A1(rf_rdata_a_ecc_i_31_), .A2(n5274), .ZN(n5636) );
NAND2_X1 U23284 ( .A1(n9294), .A2(n9295), .ZN(n768) );
NAND2_X1 U23285 ( .A1(n20947), .A2(crash_dump_o_118_), .ZN(n9295) );
NOR2_X1 U23286 ( .A1(n9296), .A2(n9297), .ZN(n9294) );
NOR2_X1 U23287 ( .A1(n11052), .A2(n8600), .ZN(n9297) );
NAND2_X1 U23288 ( .A1(n9379), .A2(n9380), .ZN(n845) );
NAND2_X1 U23289 ( .A1(n20947), .A2(crash_dump_o_116_), .ZN(n9380) );
NOR2_X1 U23290 ( .A1(n9381), .A2(n9382), .ZN(n9379) );
NOR2_X1 U23291 ( .A1(n11050), .A2(n16365), .ZN(n9382) );
NAND2_X1 U23292 ( .A1(n9465), .A2(n9466), .ZN(n926) );
NAND2_X1 U23293 ( .A1(n20947), .A2(crash_dump_o_115_), .ZN(n9466) );
NOR2_X1 U23294 ( .A1(n9467), .A2(n9468), .ZN(n9465) );
NOR2_X1 U23295 ( .A1(n11049), .A2(n16365), .ZN(n9468) );
NAND2_X1 U23296 ( .A1(n9506), .A2(n9507), .ZN(n965) );
NAND2_X1 U23297 ( .A1(n20947), .A2(crash_dump_o_114_), .ZN(n9507) );
NOR2_X1 U23298 ( .A1(n9508), .A2(n9509), .ZN(n9506) );
NOR2_X1 U23299 ( .A1(n11048), .A2(n8600), .ZN(n9509) );
NAND2_X1 U23300 ( .A1(n9550), .A2(n9551), .ZN(n1003) );
NAND2_X1 U23301 ( .A1(n20947), .A2(crash_dump_o_113_), .ZN(n9551) );
NOR2_X1 U23302 ( .A1(n9552), .A2(n9553), .ZN(n9550) );
NOR2_X1 U23303 ( .A1(n11047), .A2(n8600), .ZN(n9553) );
NAND2_X1 U23304 ( .A1(n9337), .A2(n9338), .ZN(n806) );
NAND2_X1 U23305 ( .A1(n16366), .A2(crash_dump_o_53_), .ZN(n9338) );
NOR2_X1 U23306 ( .A1(n9339), .A2(n9340), .ZN(n9337) );
NOR2_X1 U23307 ( .A1(n11495), .A2(n8773), .ZN(n9340) );
INV_X1 U23308 ( .A(rf_rdata_b_ecc_i_21_), .ZN(n20794) );
INV_X1 U23309 ( .A(rf_rdata_b_ecc_i_20_), .ZN(n20797) );
INV_X1 U23310 ( .A(rf_rdata_b_ecc_i_19_), .ZN(n20800) );
INV_X1 U23311 ( .A(rf_rdata_b_ecc_i_18_), .ZN(n20803) );
INV_X1 U23312 ( .A(rf_rdata_b_ecc_i_17_), .ZN(n20806) );
INV_X1 U23313 ( .A(rf_rdata_b_ecc_i_16_), .ZN(n20809) );
NAND2_X1 U23314 ( .A1(n6115), .A2(n6116), .ZN(n1005) );
NOR2_X1 U23315 ( .A1(n6077), .A2(n6117), .ZN(n6115) );
NAND2_X1 U23316 ( .A1(rf_rdata_b_ecc_i_17_), .A2(n20950), .ZN(n6116) );
NOR2_X1 U23317 ( .A1(n6079), .A2(n15889), .ZN(n6117) );
NAND2_X1 U23318 ( .A1(n6101), .A2(n6102), .ZN(n967) );
NOR2_X1 U23319 ( .A1(n6077), .A2(n6103), .ZN(n6101) );
NAND2_X1 U23320 ( .A1(rf_rdata_b_ecc_i_18_), .A2(n16356), .ZN(n6102) );
NOR2_X1 U23321 ( .A1(n6079), .A2(n15806), .ZN(n6103) );
NAND2_X1 U23322 ( .A1(n6075), .A2(n6076), .ZN(n928) );
NOR2_X1 U23323 ( .A1(n6077), .A2(n6078), .ZN(n6075) );
NAND2_X1 U23324 ( .A1(rf_rdata_b_ecc_i_19_), .A2(n20950), .ZN(n6076) );
NOR2_X1 U23325 ( .A1(n6079), .A2(n15885), .ZN(n6078) );
NAND2_X1 U23326 ( .A1(n6061), .A2(n6062), .ZN(n847) );
NOR2_X1 U23327 ( .A1(n5908), .A2(n6063), .ZN(n6061) );
NAND2_X1 U23328 ( .A1(rf_rdata_b_ecc_i_20_), .A2(n16356), .ZN(n6062) );
NOR2_X1 U23329 ( .A1(n11330), .A2(n5910), .ZN(n6063) );
NAND2_X1 U23330 ( .A1(n6047), .A2(n6048), .ZN(n808) );
NOR2_X1 U23331 ( .A1(n5908), .A2(n6049), .ZN(n6047) );
NAND2_X1 U23332 ( .A1(rf_rdata_b_ecc_i_21_), .A2(n20950), .ZN(n6048) );
NOR2_X1 U23333 ( .A1(n11331), .A2(n5910), .ZN(n6049) );
NAND2_X1 U23334 ( .A1(n6033), .A2(n6034), .ZN(n770) );
NOR2_X1 U23335 ( .A1(n5908), .A2(n6035), .ZN(n6033) );
NAND2_X1 U23336 ( .A1(rf_rdata_b_ecc_i_22_), .A2(n16356), .ZN(n6034) );
NOR2_X1 U23337 ( .A1(n11323), .A2(n5910), .ZN(n6035) );
INV_X1 U23338 ( .A(rf_rdata_a_ecc_i_17_), .ZN(n20680) );
INV_X1 U23339 ( .A(rf_rdata_a_ecc_i_18_), .ZN(n20646) );
INV_X1 U23340 ( .A(rf_rdata_a_ecc_i_19_), .ZN(n20608) );
INV_X1 U23341 ( .A(rf_rdata_a_ecc_i_22_), .ZN(n20488) );
INV_X1 U23342 ( .A(rf_rdata_a_ecc_i_21_), .ZN(n20528) );
INV_X1 U23343 ( .A(rf_rdata_a_ecc_i_20_), .ZN(n20568) );
NAND2_X1 U23344 ( .A1(rf_rdata_a_ecc_i_31_), .A2(n5531), .ZN(n5104) );
NAND2_X1 U23345 ( .A1(n5273), .A2(n5532), .ZN(n5531) );
NAND2_X1 U23346 ( .A1(n3952), .A2(n3953), .ZN(n3543) );
NOR2_X1 U23347 ( .A1(n3959), .A2(n3960), .ZN(n3952) );
NOR2_X1 U23348 ( .A1(n3954), .A2(n3955), .ZN(n3953) );
NOR2_X1 U23349 ( .A1(n10771), .A2(n16355), .ZN(n3960) );
NAND2_X1 U23350 ( .A1(n3941), .A2(n3942), .ZN(n3538) );
NOR2_X1 U23351 ( .A1(n3948), .A2(n3949), .ZN(n3941) );
NOR2_X1 U23352 ( .A1(n3943), .A2(n3944), .ZN(n3942) );
NOR2_X1 U23353 ( .A1(n10796), .A2(n16355), .ZN(n3949) );
NAND2_X1 U23354 ( .A1(n1865), .A2(n1866), .ZN(instr_addr_o_12_) );
NAND2_X1 U23355 ( .A1(n15929), .A2(n15991), .ZN(n1866) );
NOR2_X1 U23356 ( .A1(n1868), .A2(n1869), .ZN(n1865) );
NOR2_X1 U23357 ( .A1(n10588), .A2(n16459), .ZN(n1869) );
NAND2_X1 U23358 ( .A1(n1859), .A2(n1860), .ZN(instr_addr_o_13_) );
NAND2_X1 U23359 ( .A1(n15929), .A2(n15992), .ZN(n1860) );
NOR2_X1 U23360 ( .A1(n1862), .A2(n1863), .ZN(n1859) );
NOR2_X1 U23361 ( .A1(n10586), .A2(n16459), .ZN(n1863) );
NAND2_X1 U23362 ( .A1(n1853), .A2(n1854), .ZN(instr_addr_o_14_) );
NAND2_X1 U23363 ( .A1(n15929), .A2(n15993), .ZN(n1854) );
NOR2_X1 U23364 ( .A1(n1856), .A2(n1857), .ZN(n1853) );
NOR2_X1 U23365 ( .A1(n10584), .A2(n16459), .ZN(n1857) );
NAND2_X1 U23366 ( .A1(n1847), .A2(n1848), .ZN(instr_addr_o_15_) );
NAND2_X1 U23367 ( .A1(n15929), .A2(n15994), .ZN(n1848) );
NOR2_X1 U23368 ( .A1(n1850), .A2(n1851), .ZN(n1847) );
NOR2_X1 U23369 ( .A1(n10582), .A2(n16459), .ZN(n1851) );
INV_X1 U23370 ( .A(n23472), .ZN(n20171) );
INV_X1 U23371 ( .A(n23780), .ZN(n20109) );
INV_X1 U23372 ( .A(n23940), .ZN(n20106) );
INV_X1 U23373 ( .A(n24788), .ZN(n20334) );
INV_X1 U23374 ( .A(n24873), .ZN(n20295) );
INV_X1 U23375 ( .A(n24946), .ZN(n20256) );
INV_X1 U23376 ( .A(n24099), .ZN(n20105) );
INV_X1 U23377 ( .A(n24115), .ZN(n20162) );
INV_X1 U23378 ( .A(n24247), .ZN(n20104) );
INV_X1 U23379 ( .A(n24263), .ZN(n20160) );
INV_X1 U23380 ( .A(n24270), .ZN(n20196) );
INV_X1 U23381 ( .A(n24382), .ZN(n20103) );
INV_X1 U23382 ( .A(n24399), .ZN(n20158) );
INV_X1 U23383 ( .A(n24408), .ZN(n20194) );
INV_X1 U23384 ( .A(n24509), .ZN(n20101) );
INV_X1 U23385 ( .A(n24531), .ZN(n20156) );
INV_X1 U23386 ( .A(n24538), .ZN(n20192) );
INV_X1 U23387 ( .A(n24547), .ZN(n20228) );
INV_X1 U23388 ( .A(n24554), .ZN(n20264) );
INV_X1 U23389 ( .A(n24628), .ZN(n20100) );
INV_X1 U23390 ( .A(n24645), .ZN(n20154) );
INV_X1 U23391 ( .A(n24654), .ZN(n20190) );
INV_X1 U23392 ( .A(n24661), .ZN(n20226) );
INV_X1 U23393 ( .A(n24670), .ZN(n20262) );
INV_X1 U23394 ( .A(n24733), .ZN(n20098) );
INV_X1 U23395 ( .A(n24749), .ZN(n20152) );
INV_X1 U23396 ( .A(n24756), .ZN(n20188) );
INV_X1 U23397 ( .A(n24765), .ZN(n20224) );
INV_X1 U23398 ( .A(n24772), .ZN(n20260) );
INV_X1 U23399 ( .A(n24781), .ZN(n20297) );
INV_X1 U23400 ( .A(n24850), .ZN(n20186) );
INV_X1 U23401 ( .A(n24857), .ZN(n20222) );
INV_X1 U23402 ( .A(n24866), .ZN(n20258) );
INV_X1 U23403 ( .A(n24939), .ZN(n20220) );
NAND2_X1 U23404 ( .A1(n3930), .A2(n3931), .ZN(n3533) );
NOR2_X1 U23405 ( .A1(n3937), .A2(n3938), .ZN(n3930) );
NOR2_X1 U23406 ( .A1(n3932), .A2(n3933), .ZN(n3931) );
NOR2_X1 U23407 ( .A1(n10810), .A2(n16355), .ZN(n3938) );
NAND2_X1 U23408 ( .A1(n3919), .A2(n3920), .ZN(n3528) );
NOR2_X1 U23409 ( .A1(n3926), .A2(n3927), .ZN(n3919) );
NOR2_X1 U23410 ( .A1(n3921), .A2(n3922), .ZN(n3920) );
NOR2_X1 U23411 ( .A1(n10825), .A2(n16355), .ZN(n3927) );
NAND2_X1 U23412 ( .A1(n3896), .A2(n3897), .ZN(n3518) );
NOR2_X1 U23413 ( .A1(n3903), .A2(n3904), .ZN(n3896) );
NOR2_X1 U23414 ( .A1(n3898), .A2(n3899), .ZN(n3897) );
NOR2_X1 U23415 ( .A1(n10649), .A2(n16355), .ZN(n3904) );
INV_X1 U23416 ( .A(n24798), .ZN(n20371) );
INV_X1 U23417 ( .A(n24883), .ZN(n20332) );
INV_X1 U23418 ( .A(n24956), .ZN(n20293) );
INV_X1 U23419 ( .A(n25061), .ZN(n20215) );
INV_X1 U23420 ( .A(n25102), .ZN(n20177) );
INV_X1 U23421 ( .A(n25149), .ZN(n20139) );
INV_X1 U23422 ( .A(n25192), .ZN(n20081) );
INV_X1 U23423 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_9), .ZN(n20357) );
INV_X1 U23424 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_10), .ZN(n20320) );
INV_X1 U23425 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_11), .ZN(n20283) );
INV_X1 U23426 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_12), .ZN(n20245) );
INV_X1 U23427 ( .A(n25181), .ZN(n20029) );
INV_X1 U23428 ( .A(n25180), .ZN(n20031) );
INV_X1 U23429 ( .A(n25159), .ZN(n20087) );
INV_X1 U23430 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N45), .ZN(n20321) );
INV_X1 U23431 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N47), .ZN(n20246) );
INV_X1 U23432 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N46), .ZN(n20284) );
INV_X1 U23433 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N44), .ZN(n20358) );
INV_X1 U23434 ( .A(n25255), .ZN(n20038) );
INV_X1 U23435 ( .A(n25162), .ZN(n20035) );
INV_X1 U23436 ( .A(n25163), .ZN(n20034) );
NAND2_X1 U23437 ( .A1(n1835), .A2(n1836), .ZN(instr_addr_o_17_) );
NAND2_X1 U23438 ( .A1(n15929), .A2(n15995), .ZN(n1836) );
NOR2_X1 U23439 ( .A1(n1838), .A2(n1839), .ZN(n1835) );
NOR2_X1 U23440 ( .A1(n10578), .A2(n1706), .ZN(n1839) );
NAND2_X1 U23441 ( .A1(n1841), .A2(n1842), .ZN(instr_addr_o_16_) );
NAND2_X1 U23442 ( .A1(n15929), .A2(n16052), .ZN(n1842) );
NOR2_X1 U23443 ( .A1(n1844), .A2(n1845), .ZN(n1841) );
NOR2_X1 U23444 ( .A1(n10580), .A2(n1706), .ZN(n1845) );
NAND2_X1 U23445 ( .A1(n9089), .A2(n9090), .ZN(n575) );
NAND2_X1 U23446 ( .A1(n20947), .A2(crash_dump_o_123_), .ZN(n9090) );
NOR2_X1 U23447 ( .A1(n9091), .A2(n9092), .ZN(n9089) );
NOR2_X1 U23448 ( .A1(n11057), .A2(n16365), .ZN(n9092) );
NAND2_X1 U23449 ( .A1(n9130), .A2(n9131), .ZN(n615) );
NAND2_X1 U23450 ( .A1(n20947), .A2(crash_dump_o_122_), .ZN(n9131) );
NOR2_X1 U23451 ( .A1(n9132), .A2(n9133), .ZN(n9130) );
NOR2_X1 U23452 ( .A1(n11056), .A2(n16365), .ZN(n9133) );
NAND2_X1 U23453 ( .A1(n9171), .A2(n9172), .ZN(n655) );
NAND2_X1 U23454 ( .A1(n20947), .A2(crash_dump_o_121_), .ZN(n9172) );
NOR2_X1 U23455 ( .A1(n9173), .A2(n9174), .ZN(n9171) );
NOR2_X1 U23456 ( .A1(n11055), .A2(n8600), .ZN(n9174) );
NAND2_X1 U23457 ( .A1(n9212), .A2(n9213), .ZN(n693) );
NAND2_X1 U23458 ( .A1(n20947), .A2(crash_dump_o_120_), .ZN(n9213) );
NOR2_X1 U23459 ( .A1(n9214), .A2(n9215), .ZN(n9212) );
NOR2_X1 U23460 ( .A1(n11054), .A2(n16365), .ZN(n9215) );
NAND2_X1 U23461 ( .A1(n9253), .A2(n9254), .ZN(n730) );
NAND2_X1 U23462 ( .A1(n20947), .A2(crash_dump_o_119_), .ZN(n9254) );
NOR2_X1 U23463 ( .A1(n9255), .A2(n9256), .ZN(n9253) );
NOR2_X1 U23464 ( .A1(n11053), .A2(n8600), .ZN(n9256) );
NAND2_X1 U23465 ( .A1(n9048), .A2(n9049), .ZN(n535) );
NAND2_X1 U23466 ( .A1(n20947), .A2(crash_dump_o_124_), .ZN(n9049) );
NOR2_X1 U23467 ( .A1(n9050), .A2(n9051), .ZN(n9048) );
NOR2_X1 U23468 ( .A1(n11058), .A2(n16365), .ZN(n9051) );
INV_X1 U23469 ( .A(rf_rdata_b_ecc_i_27_), .ZN(n20776) );
INV_X1 U23470 ( .A(rf_rdata_b_ecc_i_26_), .ZN(n20779) );
INV_X1 U23471 ( .A(rf_rdata_b_ecc_i_25_), .ZN(n20782) );
INV_X1 U23472 ( .A(rf_rdata_b_ecc_i_24_), .ZN(n20785) );
INV_X1 U23473 ( .A(rf_rdata_b_ecc_i_23_), .ZN(n20788) );
INV_X1 U23474 ( .A(rf_rdata_b_ecc_i_22_), .ZN(n20791) );
NAND2_X1 U23475 ( .A1(n6019), .A2(n6020), .ZN(n732) );
NOR2_X1 U23476 ( .A1(n5908), .A2(n6021), .ZN(n6019) );
NAND2_X1 U23477 ( .A1(rf_rdata_b_ecc_i_23_), .A2(n16356), .ZN(n6020) );
NOR2_X1 U23478 ( .A1(n11332), .A2(n5910), .ZN(n6021) );
NAND2_X1 U23479 ( .A1(n6005), .A2(n6006), .ZN(n695) );
NOR2_X1 U23480 ( .A1(n5908), .A2(n6007), .ZN(n6005) );
NAND2_X1 U23481 ( .A1(rf_rdata_b_ecc_i_24_), .A2(n16356), .ZN(n6006) );
NOR2_X1 U23482 ( .A1(n11311), .A2(n5910), .ZN(n6007) );
NAND2_X1 U23483 ( .A1(n5991), .A2(n5992), .ZN(n657) );
NOR2_X1 U23484 ( .A1(n5908), .A2(n5993), .ZN(n5991) );
NAND2_X1 U23485 ( .A1(rf_rdata_b_ecc_i_25_), .A2(n16356), .ZN(n5992) );
NOR2_X1 U23486 ( .A1(n11325), .A2(n5910), .ZN(n5993) );
NAND2_X1 U23487 ( .A1(n5977), .A2(n5978), .ZN(n617) );
NOR2_X1 U23488 ( .A1(n5908), .A2(n5979), .ZN(n5977) );
NAND2_X1 U23489 ( .A1(rf_rdata_b_ecc_i_26_), .A2(n16356), .ZN(n5978) );
NOR2_X1 U23490 ( .A1(n11334), .A2(n5910), .ZN(n5979) );
NAND2_X1 U23491 ( .A1(n5963), .A2(n5964), .ZN(n577) );
NOR2_X1 U23492 ( .A1(n5908), .A2(n5965), .ZN(n5963) );
NAND2_X1 U23493 ( .A1(rf_rdata_b_ecc_i_27_), .A2(n16356), .ZN(n5964) );
NOR2_X1 U23494 ( .A1(n11336), .A2(n5910), .ZN(n5965) );
NAND2_X1 U23495 ( .A1(n5949), .A2(n5950), .ZN(n537) );
NOR2_X1 U23496 ( .A1(n5908), .A2(n5951), .ZN(n5949) );
NAND2_X1 U23497 ( .A1(rf_rdata_b_ecc_i_28_), .A2(n16356), .ZN(n5950) );
NOR2_X1 U23498 ( .A1(n11338), .A2(n5910), .ZN(n5951) );
NAND2_X1 U23499 ( .A1(n11498), .A2(n10332), .ZN(n5127) );
NAND2_X1 U23500 ( .A1(n10333), .A2(n5128), .ZN(n10332) );
NAND2_X1 U23501 ( .A1(n10334), .A2(irq_pending_o), .ZN(n10333) );
NOR2_X1 U23502 ( .A1(nmi_mode), .A2(n11477), .ZN(n10334) );
INV_X1 U23503 ( .A(rf_rdata_a_ecc_i_25_), .ZN(n20369) );
INV_X1 U23504 ( .A(rf_rdata_a_ecc_i_28_), .ZN(n20252) );
INV_X1 U23505 ( .A(rf_rdata_a_ecc_i_27_), .ZN(n20291) );
INV_X1 U23506 ( .A(rf_rdata_a_ecc_i_26_), .ZN(n20330) );
INV_X1 U23507 ( .A(rf_rdata_a_ecc_i_24_), .ZN(n20408) );
INV_X1 U23508 ( .A(rf_rdata_a_ecc_i_23_), .ZN(n20448) );
NAND2_X1 U23509 ( .A1(n10338), .A2(n10339), .ZN(n7603) );
NOR2_X1 U23510 ( .A1(n10340), .A2(n10341), .ZN(n10339) );
NOR2_X1 U23511 ( .A1(n7657), .A2(n10343), .ZN(n10338) );
NOR2_X1 U23512 ( .A1(n11483), .A2(n20892), .ZN(n10340) );
NOR2_X1 U23513 ( .A1(n11164), .A2(n20821), .ZN(n906) );
NOR2_X1 U23514 ( .A1(n11163), .A2(n20821), .ZN(n474) );
NOR2_X1 U23515 ( .A1(n11162), .A2(n20821), .ZN(n344) );
NOR2_X1 U23516 ( .A1(n11161), .A2(n20821), .ZN(n303) );
NOR2_X1 U23517 ( .A1(n11159), .A2(n20821), .ZN(n220) );
NOR2_X1 U23518 ( .A1(n11158), .A2(n20821), .ZN(n177) );
NOR2_X1 U23519 ( .A1(n11157), .A2(n20821), .ZN(n129) );
NOR2_X1 U23520 ( .A1(n11156), .A2(n20821), .ZN(n81) );
NOR2_X1 U23521 ( .A1(n11218), .A2(n20821), .ZN(n1333) );
NOR2_X1 U23522 ( .A1(n11186), .A2(n20821), .ZN(n1277) );
NOR2_X1 U23523 ( .A1(n11184), .A2(n20821), .ZN(n1238) );
NOR2_X1 U23524 ( .A1(n11183), .A2(n20821), .ZN(n1199) );
NOR2_X1 U23525 ( .A1(n11182), .A2(n20821), .ZN(n1160) );
NOR2_X1 U23526 ( .A1(n11181), .A2(n20821), .ZN(n1121) );
NAND2_X1 U23527 ( .A1(n20881), .A2(n10331), .ZN(n8056) );
NAND2_X1 U23528 ( .A1(n20991), .A2(n11517), .ZN(n10331) );
NAND2_X1 U23529 ( .A1(n3997), .A2(n3998), .ZN(n3402) );
NOR2_X1 U23530 ( .A1(n4007), .A2(n4008), .ZN(n3997) );
NOR2_X1 U23531 ( .A1(n3999), .A2(n4000), .ZN(n3998) );
NOR2_X1 U23532 ( .A1(n10730), .A2(n20931), .ZN(n4008) );
NAND2_X1 U23533 ( .A1(n3986), .A2(n3987), .ZN(n3397) );
NOR2_X1 U23534 ( .A1(n3993), .A2(n3994), .ZN(n3986) );
NOR2_X1 U23535 ( .A1(n3988), .A2(n3989), .ZN(n3987) );
NOR2_X1 U23536 ( .A1(n10744), .A2(n16355), .ZN(n3994) );
NAND2_X1 U23537 ( .A1(n1877), .A2(n1878), .ZN(instr_addr_o_10_) );
NAND2_X1 U23538 ( .A1(n15929), .A2(n15996), .ZN(n1878) );
NOR2_X1 U23539 ( .A1(n1880), .A2(n1881), .ZN(n1877) );
NOR2_X1 U23540 ( .A1(n10592), .A2(n16459), .ZN(n1881) );
NAND2_X1 U23541 ( .A1(n1871), .A2(n1872), .ZN(instr_addr_o_11_) );
NAND2_X1 U23542 ( .A1(n15929), .A2(n16051), .ZN(n1872) );
NOR2_X1 U23543 ( .A1(n1874), .A2(n1875), .ZN(n1871) );
NOR2_X1 U23544 ( .A1(n10590), .A2(n16459), .ZN(n1875) );
NAND2_X1 U23545 ( .A1(n1721), .A2(n1722), .ZN(instr_addr_o_6_) );
NAND2_X1 U23546 ( .A1(n15929), .A2(n15997), .ZN(n1722) );
NOR2_X1 U23547 ( .A1(n1724), .A2(n1725), .ZN(n1721) );
NOR2_X1 U23548 ( .A1(n10600), .A2(n16459), .ZN(n1725) );
NAND2_X1 U23549 ( .A1(n1709), .A2(n1710), .ZN(instr_addr_o_8_) );
NAND2_X1 U23550 ( .A1(n15929), .A2(n15998), .ZN(n1710) );
NOR2_X1 U23551 ( .A1(n1712), .A2(n1713), .ZN(n1709) );
NOR2_X1 U23552 ( .A1(n10596), .A2(n16459), .ZN(n1713) );
NAND2_X1 U23553 ( .A1(n1700), .A2(n1701), .ZN(instr_addr_o_9_) );
NAND2_X1 U23554 ( .A1(n15929), .A2(n15999), .ZN(n1701) );
NOR2_X1 U23555 ( .A1(n1704), .A2(n1705), .ZN(n1700) );
NOR2_X1 U23556 ( .A1(n10594), .A2(n16459), .ZN(n1705) );
NOR2_X1 U23557 ( .A1(n261), .A2(n262), .ZN(n258) );
NOR2_X1 U23558 ( .A1(n83), .A2(n16241), .ZN(n261) );
NOR2_X1 U23559 ( .A1(n11160), .A2(n20821), .ZN(n262) );
INV_X1 U23560 ( .A(n25009), .ZN(n20218) );
INV_X1 U23561 ( .A(n25060), .ZN(n20180) );
INV_X1 U23562 ( .A(n25101), .ZN(n20142) );
INV_X1 U23563 ( .A(n24824), .ZN(n20097) );
INV_X1 U23564 ( .A(n24841), .ZN(n20150) );
INV_X1 U23565 ( .A(n24907), .ZN(n20095) );
INV_X1 U23566 ( .A(n24923), .ZN(n20148) );
INV_X1 U23567 ( .A(n24930), .ZN(n20184) );
INV_X1 U23568 ( .A(n24976), .ZN(n20094) );
INV_X1 U23569 ( .A(n24993), .ZN(n20146) );
INV_X1 U23570 ( .A(n25002), .ZN(n20182) );
INV_X1 U23571 ( .A(n25037), .ZN(n20092) );
INV_X1 U23572 ( .A(n25053), .ZN(n20144) );
INV_X1 U23573 ( .A(n25084), .ZN(n20091) );
INV_X1 U23574 ( .A(n25123), .ZN(n20089) );
NAND2_X1 U23575 ( .A1(n10335), .A2(n7628), .ZN(irq_pending_o) );
NOR2_X1 U23576 ( .A1(n10337), .A2(n7603), .ZN(n10335) );
NOR2_X1 U23577 ( .A1(n11309), .A2(n20882), .ZN(n10337) );
NAND2_X1 U23578 ( .A1(n10314), .A2(n16439), .ZN(n3703) );
NOR2_X1 U23579 ( .A1(n11459), .A2(n10460), .ZN(n10314) );
NOR2_X1 U23580 ( .A1(n15927), .A2(n15812), .ZN(n10460) );
NAND2_X1 U23581 ( .A1(irq_fast_i_9_), .A2(n16000), .ZN(n7654) );
NAND2_X1 U23582 ( .A1(irq_fast_i_10_), .A2(n16001), .ZN(n7693) );
NAND2_X1 U23583 ( .A1(n4011), .A2(n4012), .ZN(n3407) );
NOR2_X1 U23584 ( .A1(n4014), .A2(n4015), .ZN(n4011) );
NOR2_X1 U23585 ( .A1(n16428), .A2(n4013), .ZN(n4012) );
NOR2_X1 U23586 ( .A1(n10682), .A2(n16355), .ZN(n4015) );
NAND2_X1 U23587 ( .A1(n4018), .A2(n4019), .ZN(n3412) );
NOR2_X1 U23588 ( .A1(n4022), .A2(n4023), .ZN(n4018) );
NOR2_X1 U23589 ( .A1(n4020), .A2(n4021), .ZN(n4019) );
NOR2_X1 U23590 ( .A1(n10716), .A2(n20931), .ZN(n4023) );
NAND2_X1 U23591 ( .A1(n3975), .A2(n3976), .ZN(n3553) );
NOR2_X1 U23592 ( .A1(n3982), .A2(n3983), .ZN(n3975) );
NOR2_X1 U23593 ( .A1(n3977), .A2(n3978), .ZN(n3976) );
NOR2_X1 U23594 ( .A1(n10758), .A2(n16355), .ZN(n3983) );
INV_X1 U23595 ( .A(n25019), .ZN(n20254) );
INV_X1 U23596 ( .A(n25070), .ZN(n20216) );
INV_X1 U23597 ( .A(n25111), .ZN(n20178) );
INV_X1 U23598 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_5), .ZN(n20507) );
INV_X1 U23599 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_6), .ZN(n20469) );
INV_X1 U23600 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_7), .ZN(n20431) );
INV_X1 U23601 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_8), .ZN(n20394) );
NAND2_X1 U23602 ( .A1(n9979), .A2(n9980), .ZN(n9978) );
NAND2_X1 U23603 ( .A1(n9987), .A2(n197), .ZN(n9979) );
NAND2_X1 U23604 ( .A1(n11498), .A2(n9981), .ZN(n9980) );
NAND2_X1 U23605 ( .A1(n9988), .A2(n9989), .ZN(n9987) );
INV_X1 U23606 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N41), .ZN(n20470) );
INV_X1 U23607 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N43), .ZN(n20395) );
INV_X1 U23608 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N40), .ZN(n20508) );
INV_X1 U23609 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N42), .ZN(n20432) );
NAND2_X1 U23610 ( .A1(n11471), .A2(n10311), .ZN(instr_req_o) );
NAND2_X1 U23611 ( .A1(n10312), .A2(n10313), .ZN(n10311) );
NOR2_X1 U23612 ( .A1(n20895), .A2(n15878), .ZN(n10312) );
AND2_X1 U23613 ( .A1(n3704), .A2(n3703), .ZN(n10313) );
NAND2_X1 U23614 ( .A1(n1715), .A2(n1716), .ZN(instr_addr_o_7_) );
NAND2_X1 U23615 ( .A1(n15929), .A2(n16002), .ZN(n1716) );
NOR2_X1 U23616 ( .A1(n1718), .A2(n1719), .ZN(n1715) );
NOR2_X1 U23617 ( .A1(n10598), .A2(n16459), .ZN(n1719) );
NAND2_X1 U23618 ( .A1(n8962), .A2(n8963), .ZN(n414) );
NAND2_X1 U23619 ( .A1(n16366), .A2(crash_dump_o_62_), .ZN(n8963) );
NOR2_X1 U23620 ( .A1(n8964), .A2(n8965), .ZN(n8962) );
NOR2_X1 U23621 ( .A1(n11505), .A2(n8773), .ZN(n8965) );
NAND2_X1 U23622 ( .A1(n10131), .A2(n10132), .ZN(n5799) );
NAND2_X1 U23623 ( .A1(n16366), .A2(crash_dump_o_63_), .ZN(n10132) );
NOR2_X1 U23624 ( .A1(n10135), .A2(n10136), .ZN(n10131) );
NOR2_X1 U23625 ( .A1(n11467), .A2(n8773), .ZN(n10136) );
NAND2_X1 U23626 ( .A1(n9007), .A2(n9008), .ZN(n495) );
NAND2_X1 U23627 ( .A1(n20947), .A2(crash_dump_o_125_), .ZN(n9008) );
NOR2_X1 U23628 ( .A1(n9009), .A2(n9010), .ZN(n9007) );
NOR2_X1 U23629 ( .A1(n11492), .A2(n16365), .ZN(n9010) );
INV_X1 U23630 ( .A(rf_rdata_b_ecc_i_30_), .ZN(n20767) );
INV_X1 U23631 ( .A(rf_rdata_b_ecc_i_29_), .ZN(n20770) );
INV_X1 U23632 ( .A(rf_rdata_b_ecc_i_28_), .ZN(n20773) );
NAND2_X1 U23633 ( .A1(n5925), .A2(n5926), .ZN(n497) );
NOR2_X1 U23634 ( .A1(n5908), .A2(n5927), .ZN(n5925) );
NAND2_X1 U23635 ( .A1(rf_rdata_b_ecc_i_29_), .A2(n16356), .ZN(n5926) );
NOR2_X1 U23636 ( .A1(n11493), .A2(n5910), .ZN(n5927) );
NOR2_X1 U23637 ( .A1(n10772), .A2(n8575), .ZN(n9724) );
NOR2_X1 U23638 ( .A1(n10761), .A2(n8575), .ZN(n9763) );
NOR2_X1 U23639 ( .A1(n10720), .A2(n8575), .ZN(n8616) );
NOR2_X1 U23640 ( .A1(n10684), .A2(n8575), .ZN(n8659) );
NOR2_X1 U23641 ( .A1(n10665), .A2(n8575), .ZN(n9904) );
NOR2_X1 U23642 ( .A1(n10667), .A2(n8575), .ZN(n9858) );
NOR2_X1 U23643 ( .A1(n10666), .A2(n8575), .ZN(n9398) );
NOR2_X1 U23644 ( .A1(n11114), .A2(n8575), .ZN(n9312) );
NOR2_X1 U23645 ( .A1(n10650), .A2(n8575), .ZN(n9524) );
NOR2_X1 U23646 ( .A1(n10873), .A2(n8575), .ZN(n9356) );
NOR2_X1 U23647 ( .A1(n10811), .A2(n8575), .ZN(n9617) );
NOR2_X1 U23648 ( .A1(n10797), .A2(n8575), .ZN(n9654) );
NOR2_X1 U23649 ( .A1(n10782), .A2(n8575), .ZN(n9691) );
NOR2_X1 U23650 ( .A1(n10747), .A2(n8575), .ZN(n9816) );
NOR2_X1 U23651 ( .A1(n10734), .A2(n8575), .ZN(n8574) );
NOR2_X1 U23652 ( .A1(n10707), .A2(n8575), .ZN(n8713) );
NOR2_X1 U23653 ( .A1(n11115), .A2(n8575), .ZN(n8939) );
NOR2_X1 U23654 ( .A1(n10976), .A2(n8685), .ZN(n9085) );
NOR2_X1 U23655 ( .A1(n10961), .A2(n8685), .ZN(n9126) );
NOR2_X1 U23656 ( .A1(n10946), .A2(n8685), .ZN(n9167) );
NOR2_X1 U23657 ( .A1(n10931), .A2(n8685), .ZN(n9208) );
NOR2_X1 U23658 ( .A1(n10916), .A2(n8685), .ZN(n9249) );
NOR2_X1 U23659 ( .A1(n10901), .A2(n8685), .ZN(n9290) );
NOR2_X1 U23660 ( .A1(n10871), .A2(n8685), .ZN(n9461) );
NOR2_X1 U23661 ( .A1(n10856), .A2(n8685), .ZN(n9502) );
NOR2_X1 U23662 ( .A1(n10839), .A2(n8685), .ZN(n9588) );
NOR2_X1 U23663 ( .A1(n11489), .A2(n8685), .ZN(n9044) );
NOR2_X1 U23664 ( .A1(n11147), .A2(n8685), .ZN(n9003) );
NAND2_X1 U23665 ( .A1(irq_nm_i), .A2(n15919), .ZN(n5128) );
NOR2_X1 U23666 ( .A1(n10995), .A2(n16368), .ZN(n9364) );
NOR2_X1 U23667 ( .A1(n10988), .A2(n16368), .ZN(n9087) );
NOR2_X1 U23668 ( .A1(n10989), .A2(n16368), .ZN(n9128) );
NOR2_X1 U23669 ( .A1(n10990), .A2(n16368), .ZN(n9169) );
NOR2_X1 U23670 ( .A1(n10991), .A2(n16368), .ZN(n9210) );
NOR2_X1 U23671 ( .A1(n10992), .A2(n16368), .ZN(n9251) );
NOR2_X1 U23672 ( .A1(n10993), .A2(n16368), .ZN(n9292) );
NOR2_X1 U23673 ( .A1(n10996), .A2(n16367), .ZN(n9463) );
NOR2_X1 U23674 ( .A1(n10997), .A2(n16367), .ZN(n9504) );
NOR2_X1 U23675 ( .A1(n10999), .A2(n16367), .ZN(n9590) );
NOR2_X1 U23676 ( .A1(n10820), .A2(n16367), .ZN(n9628) );
NOR2_X1 U23677 ( .A1(n11000), .A2(n16367), .ZN(n9665) );
NOR2_X1 U23678 ( .A1(n10791), .A2(n16367), .ZN(n9702) );
NOR2_X1 U23679 ( .A1(n11302), .A2(n16367), .ZN(n9722) );
NOR2_X1 U23680 ( .A1(n11001), .A2(n16367), .ZN(n9772) );
NOR2_X1 U23681 ( .A1(n11002), .A2(n16367), .ZN(n9827) );
NOR2_X1 U23682 ( .A1(n11003), .A2(n16367), .ZN(n8592) );
NOR2_X1 U23683 ( .A1(n11303), .A2(n16368), .ZN(n9934) );
NOR2_X1 U23684 ( .A1(n11301), .A2(n16367), .ZN(n9875) );
NOR2_X1 U23685 ( .A1(n10780), .A2(n16368), .ZN(n9412) );
NOR2_X1 U23686 ( .A1(n10987), .A2(n16368), .ZN(n9046) );
NOR2_X1 U23687 ( .A1(n10986), .A2(n16368), .ZN(n9005) );
NOR2_X1 U23688 ( .A1(n10994), .A2(n16368), .ZN(n9321) );
NOR2_X1 U23689 ( .A1(n10998), .A2(n16367), .ZN(n9533) );
NOR2_X1 U23690 ( .A1(n10794), .A2(n16385), .ZN(n9686) );
NOR2_X1 U23691 ( .A1(n10756), .A2(n16385), .ZN(n9811) );
NOR2_X1 U23692 ( .A1(n10823), .A2(n16385), .ZN(n9612) );
NOR2_X1 U23693 ( .A1(n10808), .A2(n16385), .ZN(n9649) );
INV_X1 U23694 ( .A(rf_rdata_a_ecc_i_29_), .ZN(n20214) );
INV_X1 U23695 ( .A(rf_rdata_a_ecc_i_31_), .ZN(n20137) );
INV_X1 U23696 ( .A(rf_rdata_a_ecc_i_30_), .ZN(n20176) );
NOR2_X1 U23697 ( .A1(n11103), .A2(n8102), .ZN(n9928) );
NOR2_X1 U23698 ( .A1(n11112), .A2(n8102), .ZN(n9869) );
NOR2_X1 U23699 ( .A1(n11113), .A2(n16385), .ZN(n9406) );
NOR2_X1 U23700 ( .A1(n10733), .A2(n8576), .ZN(n8573) );
NOR2_X1 U23701 ( .A1(n10743), .A2(n16369), .ZN(n8588) );
NOR2_X1 U23702 ( .A1(n10729), .A2(n16369), .ZN(n8633) );
NOR2_X1 U23703 ( .A1(n10706), .A2(n8576), .ZN(n8712) );
NOR2_X1 U23704 ( .A1(n10715), .A2(n16369), .ZN(n8722) );
NOR2_X1 U23705 ( .A1(n10699), .A2(n8585), .ZN(n8804) );
NOR2_X1 U23706 ( .A1(n10702), .A2(n16369), .ZN(n8809) );
NOR2_X1 U23707 ( .A1(n10693), .A2(n8576), .ZN(n8795) );
NOR2_X1 U23708 ( .A1(n10679), .A2(n16372), .ZN(n8679) );
NOR2_X1 U23709 ( .A1(n10675), .A2(n16375), .ZN(n8835) );
NOR2_X1 U23710 ( .A1(n10981), .A2(n16372), .ZN(n8915) );
NOR2_X1 U23711 ( .A1(n10618), .A2(n8585), .ZN(n8919) );
NOR2_X1 U23712 ( .A1(n11134), .A2(n16369), .ZN(n8921) );
NOR2_X1 U23713 ( .A1(n10613), .A2(n8576), .ZN(n8906) );
NOR2_X1 U23714 ( .A1(n11016), .A2(n8585), .ZN(n8764) );
NOR2_X1 U23715 ( .A1(n11119), .A2(n8576), .ZN(n8749) );
NOR2_X1 U23716 ( .A1(n10722), .A2(n16375), .ZN(n8617) );
NOR2_X1 U23717 ( .A1(n10719), .A2(n8576), .ZN(n8619) );
NOR2_X1 U23718 ( .A1(n10726), .A2(n8585), .ZN(n8636) );
NOR2_X1 U23719 ( .A1(n10686), .A2(n16375), .ZN(n8660) );
NOR2_X1 U23720 ( .A1(n10683), .A2(n8576), .ZN(n8662) );
NOR2_X1 U23721 ( .A1(n10687), .A2(n8585), .ZN(n8676) );
NOR2_X1 U23722 ( .A1(n10673), .A2(n8576), .ZN(n8840) );
NOR2_X1 U23723 ( .A1(n8863), .A2(n8864), .ZN(n8861) );
NOR2_X1 U23724 ( .A1(n11144), .A2(n8685), .ZN(n8863) );
NOR2_X1 U23725 ( .A1(n11141), .A2(n16369), .ZN(n8864) );
NOR2_X1 U23726 ( .A1(n11140), .A2(n16369), .ZN(n8765) );
NOR2_X1 U23727 ( .A1(n10610), .A2(n16372), .ZN(n8767) );
NOR2_X1 U23728 ( .A1(n10742), .A2(n16385), .ZN(n8566) );
NOR2_X1 U23729 ( .A1(n10714), .A2(n16385), .ZN(n8708) );
NAND2_X1 U23730 ( .A1(n5905), .A2(n5906), .ZN(n412) );
NOR2_X1 U23731 ( .A1(n5908), .A2(n5909), .ZN(n5905) );
NAND2_X1 U23732 ( .A1(rf_rdata_b_ecc_i_30_), .A2(n16356), .ZN(n5906) );
NOR2_X1 U23733 ( .A1(n11340), .A2(n5910), .ZN(n5909) );
NOR2_X1 U23734 ( .A1(n10983), .A2(n16368), .ZN(n8635) );
NOR2_X1 U23735 ( .A1(n10777), .A2(n16367), .ZN(n8724) );
NOR2_X1 U23736 ( .A1(n11005), .A2(n16368), .ZN(n8811) );
NOR2_X1 U23737 ( .A1(n10982), .A2(n16367), .ZN(n8669) );
NOR2_X1 U23738 ( .A1(n11006), .A2(n16368), .ZN(n8847) );
NOR2_X1 U23739 ( .A1(n10985), .A2(n16367), .ZN(n8947) );
NAND2_X1 U23740 ( .A1(irq_fast_i_6_), .A2(n16003), .ZN(n7658) );
NOR2_X1 U23741 ( .A1(n10887), .A2(n16383), .ZN(n9355) );
NOR2_X1 U23742 ( .A1(n11507), .A2(n16383), .ZN(n8938) );
NOR2_X1 U23743 ( .A1(n10612), .A2(n8806), .ZN(n8920) );
NOR2_X1 U23744 ( .A1(n10824), .A2(n8591), .ZN(n9626) );
NOR2_X1 U23745 ( .A1(n10809), .A2(n8591), .ZN(n9663) );
NOR2_X1 U23746 ( .A1(n10795), .A2(n8591), .ZN(n9700) );
NOR2_X1 U23747 ( .A1(n10979), .A2(n8584), .ZN(n9783) );
NOR2_X1 U23748 ( .A1(n10757), .A2(n8591), .ZN(n9825) );
NOR2_X1 U23749 ( .A1(n11009), .A2(n16371), .ZN(n9936) );
NOR2_X1 U23750 ( .A1(n11014), .A2(n16371), .ZN(n9877) );
NOR2_X1 U23751 ( .A1(n11012), .A2(n8585), .ZN(n9414) );
NOR2_X1 U23752 ( .A1(n10617), .A2(n8584), .ZN(n9329) );
NOR2_X1 U23753 ( .A1(n10646), .A2(n8584), .ZN(n9542) );
NOR2_X1 U23754 ( .A1(n10964), .A2(n16373), .ZN(n9072) );
NOR2_X1 U23755 ( .A1(n10949), .A2(n16373), .ZN(n9113) );
NOR2_X1 U23756 ( .A1(n10934), .A2(n16373), .ZN(n9154) );
NOR2_X1 U23757 ( .A1(n10919), .A2(n16373), .ZN(n9195) );
NOR2_X1 U23758 ( .A1(n10904), .A2(n16373), .ZN(n9236) );
NOR2_X1 U23759 ( .A1(n10889), .A2(n16373), .ZN(n9277) );
NOR2_X1 U23760 ( .A1(n10874), .A2(n16373), .ZN(n9375) );
NOR2_X1 U23761 ( .A1(n10859), .A2(n8576), .ZN(n9448) );
NOR2_X1 U23762 ( .A1(n10842), .A2(n8576), .ZN(n9489) );
NOR2_X1 U23763 ( .A1(n10827), .A2(n8576), .ZN(n9575) );
NOR2_X1 U23764 ( .A1(n10812), .A2(n8576), .ZN(n9616) );
NOR2_X1 U23765 ( .A1(n10798), .A2(n8576), .ZN(n9653) );
NOR2_X1 U23766 ( .A1(n10783), .A2(n8576), .ZN(n9690) );
NOR2_X1 U23767 ( .A1(n10775), .A2(n8572), .ZN(n9740) );
NOR2_X1 U23768 ( .A1(n10748), .A2(n8576), .ZN(n9815) );
NOR2_X1 U23769 ( .A1(n10636), .A2(n16373), .ZN(n9031) );
NOR2_X1 U23770 ( .A1(n10626), .A2(n16373), .ZN(n8990) );
NOR2_X1 U23771 ( .A1(n11508), .A2(n16373), .ZN(n8958) );
NOR2_X1 U23772 ( .A1(n10977), .A2(n16383), .ZN(n9075) );
NOR2_X1 U23773 ( .A1(n10962), .A2(n8104), .ZN(n9116) );
NOR2_X1 U23774 ( .A1(n10947), .A2(n8104), .ZN(n9157) );
NOR2_X1 U23775 ( .A1(n10932), .A2(n8104), .ZN(n9198) );
NOR2_X1 U23776 ( .A1(n10917), .A2(n8104), .ZN(n9239) );
NOR2_X1 U23777 ( .A1(n10902), .A2(n8104), .ZN(n9280) );
NOR2_X1 U23778 ( .A1(n10872), .A2(n16383), .ZN(n9451) );
NOR2_X1 U23779 ( .A1(n10857), .A2(n16383), .ZN(n9492) );
NOR2_X1 U23780 ( .A1(n10840), .A2(n16383), .ZN(n9578) );
NOR2_X1 U23781 ( .A1(n10825), .A2(n16383), .ZN(n9629) );
NOR2_X1 U23782 ( .A1(n10810), .A2(n16383), .ZN(n9666) );
NOR2_X1 U23783 ( .A1(n10796), .A2(n16383), .ZN(n9703) );
NOR2_X1 U23784 ( .A1(n11306), .A2(n16383), .ZN(n9773) );
NOR2_X1 U23785 ( .A1(n10758), .A2(n16383), .ZN(n9828) );
NOR2_X1 U23786 ( .A1(n10781), .A2(n16383), .ZN(n9935) );
NOR2_X1 U23787 ( .A1(n10664), .A2(n16383), .ZN(n9876) );
NOR2_X1 U23788 ( .A1(n11486), .A2(n16383), .ZN(n9413) );
NOR2_X1 U23789 ( .A1(n10634), .A2(n8104), .ZN(n9034) );
NOR2_X1 U23790 ( .A1(n10624), .A2(n8104), .ZN(n8993) );
NOR2_X1 U23791 ( .A1(n11497), .A2(n16383), .ZN(n9322) );
NOR2_X1 U23792 ( .A1(n10649), .A2(n16383), .ZN(n9534) );
NOR2_X1 U23793 ( .A1(n10968), .A2(n16372), .ZN(n9082) );
NOR2_X1 U23794 ( .A1(n10953), .A2(n16372), .ZN(n9123) );
NOR2_X1 U23795 ( .A1(n10938), .A2(n16372), .ZN(n9164) );
NOR2_X1 U23796 ( .A1(n10923), .A2(n16372), .ZN(n9205) );
NOR2_X1 U23797 ( .A1(n10908), .A2(n16372), .ZN(n9246) );
NOR2_X1 U23798 ( .A1(n10893), .A2(n8584), .ZN(n9287) );
NOR2_X1 U23799 ( .A1(n10882), .A2(n8585), .ZN(n9378) );
NOR2_X1 U23800 ( .A1(n10863), .A2(n8584), .ZN(n9458) );
NOR2_X1 U23801 ( .A1(n10846), .A2(n8584), .ZN(n9499) );
NOR2_X1 U23802 ( .A1(n10831), .A2(n8584), .ZN(n9585) );
NOR2_X1 U23803 ( .A1(n11010), .A2(n16371), .ZN(n9779) );
NOR2_X1 U23804 ( .A1(n10631), .A2(n16372), .ZN(n9041) );
NOR2_X1 U23805 ( .A1(n10621), .A2(n8584), .ZN(n9000) );
NOR2_X1 U23806 ( .A1(n10619), .A2(n8585), .ZN(n8961) );
NOR2_X1 U23807 ( .A1(n11013), .A2(n16371), .ZN(n9328) );
NOR2_X1 U23808 ( .A1(n10656), .A2(n16371), .ZN(n9540) );
NOR2_X1 U23809 ( .A1(n10608), .A2(n16459), .ZN(n1761) );
NOR2_X1 U23810 ( .A1(n10606), .A2(n1706), .ZN(n1743) );
NOR2_X1 U23811 ( .A1(n10604), .A2(n1706), .ZN(n1737) );
NOR2_X1 U23812 ( .A1(n10876), .A2(n16374), .ZN(n9358) );
NOR2_X1 U23813 ( .A1(n10774), .A2(n8567), .ZN(n9725) );
NOR2_X1 U23814 ( .A1(n10773), .A2(n16373), .ZN(n9741) );
NOR2_X1 U23815 ( .A1(n10763), .A2(n8567), .ZN(n9764) );
NOR2_X1 U23816 ( .A1(n10762), .A2(n16373), .ZN(n9766) );
NOR2_X1 U23817 ( .A1(n11479), .A2(n8567), .ZN(n9905) );
NOR2_X1 U23818 ( .A1(n11116), .A2(n8576), .ZN(n9912) );
NOR2_X1 U23819 ( .A1(n11124), .A2(n8567), .ZN(n9859) );
NOR2_X1 U23820 ( .A1(n11118), .A2(n8576), .ZN(n9861) );
NOR2_X1 U23821 ( .A1(n11122), .A2(n16375), .ZN(n9399) );
NOR2_X1 U23822 ( .A1(n11117), .A2(n16373), .ZN(n9401) );
NOR2_X1 U23823 ( .A1(n10628), .A2(n16374), .ZN(n8941) );
NOR2_X1 U23824 ( .A1(n11123), .A2(n16375), .ZN(n9313) );
NOR2_X1 U23825 ( .A1(n11120), .A2(n16373), .ZN(n9315) );
NOR2_X1 U23826 ( .A1(n10652), .A2(n8567), .ZN(n9525) );
NOR2_X1 U23827 ( .A1(n10651), .A2(n8576), .ZN(n9527) );
NOR2_X1 U23828 ( .A1(n10688), .A2(n16362), .ZN(n8665) );
NOR2_X1 U23829 ( .A1(n11100), .A2(n8624), .ZN(n8846) );
NOR2_X1 U23830 ( .A1(n11094), .A2(n16362), .ZN(n8946) );
NOR2_X1 U23831 ( .A1(n10883), .A2(n16362), .ZN(n9363) );
NOR2_X1 U23832 ( .A1(n11098), .A2(n16362), .ZN(n9769) );
NOR2_X1 U23833 ( .A1(n11096), .A2(n16362), .ZN(n9318) );
NOR2_X1 U23834 ( .A1(n10657), .A2(n16362), .ZN(n9530) );
NOR2_X1 U23835 ( .A1(n11480), .A2(n16361), .ZN(n9864) );
NAND2_X1 U23836 ( .A1(n5892), .A2(n5893), .ZN(n5891) );
NAND2_X1 U23837 ( .A1(n11216), .A2(n20958), .ZN(n5893) );
NAND2_X1 U23838 ( .A1(n5818), .A2(n20137), .ZN(n5892) );
NOR2_X1 U23839 ( .A1(n10973), .A2(n16362), .ZN(n9073) );
NOR2_X1 U23840 ( .A1(n10958), .A2(n16362), .ZN(n9114) );
NOR2_X1 U23841 ( .A1(n10943), .A2(n16362), .ZN(n9155) );
NOR2_X1 U23842 ( .A1(n10700), .A2(n16362), .ZN(n8798) );
NOR2_X1 U23843 ( .A1(n10640), .A2(n16362), .ZN(n9032) );
NOR2_X1 U23844 ( .A1(n11095), .A2(n16362), .ZN(n8991) );
NOR2_X1 U23845 ( .A1(n11093), .A2(n16362), .ZN(n8907) );
NOR2_X1 U23846 ( .A1(n11099), .A2(n16362), .ZN(n8753) );
NOR2_X1 U23847 ( .A1(n10928), .A2(n16362), .ZN(n9196) );
NOR2_X1 U23848 ( .A1(n10913), .A2(n16362), .ZN(n9237) );
NOR2_X1 U23849 ( .A1(n10898), .A2(n16362), .ZN(n9278) );
NOR2_X1 U23850 ( .A1(n10868), .A2(n16362), .ZN(n9449) );
NOR2_X1 U23851 ( .A1(n10851), .A2(n16362), .ZN(n9490) );
NOR2_X1 U23852 ( .A1(n10836), .A2(n16362), .ZN(n9576) );
NOR2_X1 U23853 ( .A1(n11102), .A2(n16362), .ZN(n9407) );
NOR2_X1 U23854 ( .A1(n11509), .A2(n16361), .ZN(n9922) );
NOR2_X1 U23855 ( .A1(n11310), .A2(n16361), .ZN(n9405) );
AND2_X1 U23856 ( .A1(irq_fast_i_14_), .A2(n16127), .ZN(n7643) );
NOR2_X1 U23857 ( .A1(n10779), .A2(n8688), .ZN(n9742) );
NOR2_X1 U23858 ( .A1(n11149), .A2(n8751), .ZN(n9921) );
NAND2_X1 U23859 ( .A1(n9873), .A2(n9874), .ZN(n9872) );
NOR2_X1 U23860 ( .A1(n9877), .A2(n9878), .ZN(n9873) );
NOR2_X1 U23861 ( .A1(n9875), .A2(n9876), .ZN(n9874) );
NOR2_X1 U23862 ( .A1(n11482), .A2(n8806), .ZN(n9878) );
NAND2_X1 U23863 ( .A1(n9410), .A2(n9411), .ZN(n9409) );
NOR2_X1 U23864 ( .A1(n9414), .A2(n9415), .ZN(n9410) );
NOR2_X1 U23865 ( .A1(n9412), .A2(n9413), .ZN(n9411) );
NOR2_X1 U23866 ( .A1(n11488), .A2(n8806), .ZN(n9415) );
NOR2_X1 U23867 ( .A1(n11150), .A2(n8751), .ZN(n8796) );
NOR2_X1 U23868 ( .A1(n11521), .A2(n8751), .ZN(n8750) );
NOR2_X1 U23869 ( .A1(n7679), .A2(n7657), .ZN(n7676) );
NOR2_X1 U23870 ( .A1(n7680), .A2(n7681), .ZN(n7679) );
NOR2_X1 U23871 ( .A1(n10916), .A2(n20891), .ZN(n7681) );
NOR2_X1 U23872 ( .A1(n20890), .A2(n7683), .ZN(n7680) );
NOR2_X1 U23873 ( .A1(n11293), .A2(n6541), .ZN(n6538) );
NOR2_X1 U23874 ( .A1(n6542), .A2(n1590), .ZN(n6541) );
NOR2_X1 U23875 ( .A1(n20935), .A2(n6318), .ZN(n6542) );
NOR2_X1 U23876 ( .A1(n4047), .A2(n4048), .ZN(n4044) );
NOR2_X1 U23877 ( .A1(n4054), .A2(n20983), .ZN(n4047) );
NOR2_X1 U23878 ( .A1(n3777), .A2(n4049), .ZN(n4048) );
NOR2_X1 U23879 ( .A1(n11498), .A2(n4056), .ZN(n4054) );
NOR2_X1 U23880 ( .A1(n7694), .A2(n20889), .ZN(n7690) );
NOR2_X1 U23881 ( .A1(n7696), .A2(n7697), .ZN(n7694) );
NAND2_X1 U23882 ( .A1(n7698), .A2(n7651), .ZN(n7696) );
NAND2_X1 U23883 ( .A1(n7684), .A2(irq_fast_i_1_), .ZN(n7697) );
NAND2_X1 U23884 ( .A1(n9624), .A2(n9625), .ZN(n9618) );
NOR2_X1 U23885 ( .A1(n9626), .A2(n9627), .ZN(n9625) );
NOR2_X1 U23886 ( .A1(n9628), .A2(n9629), .ZN(n9624) );
NOR2_X1 U23887 ( .A1(n10819), .A2(n8590), .ZN(n9627) );
NAND2_X1 U23888 ( .A1(n9661), .A2(n9662), .ZN(n9655) );
NOR2_X1 U23889 ( .A1(n9663), .A2(n9664), .ZN(n9662) );
NOR2_X1 U23890 ( .A1(n9665), .A2(n9666), .ZN(n9661) );
NOR2_X1 U23891 ( .A1(n10805), .A2(n8590), .ZN(n9664) );
NAND2_X1 U23892 ( .A1(n9698), .A2(n9699), .ZN(n9692) );
NOR2_X1 U23893 ( .A1(n9700), .A2(n9701), .ZN(n9699) );
NOR2_X1 U23894 ( .A1(n9702), .A2(n9703), .ZN(n9698) );
NOR2_X1 U23895 ( .A1(n10790), .A2(n8590), .ZN(n9701) );
NAND2_X1 U23896 ( .A1(n9823), .A2(n9824), .ZN(n9817) );
NOR2_X1 U23897 ( .A1(n9825), .A2(n9826), .ZN(n9824) );
NOR2_X1 U23898 ( .A1(n9827), .A2(n9828), .ZN(n9823) );
NOR2_X1 U23899 ( .A1(n10751), .A2(n8590), .ZN(n9826) );
NOR2_X1 U23900 ( .A1(n10744), .A2(n16383), .ZN(n8593) );
NOR2_X1 U23901 ( .A1(n10716), .A2(n16383), .ZN(n8725) );
NOR2_X1 U23902 ( .A1(n10703), .A2(n16383), .ZN(n8812) );
NOR2_X1 U23903 ( .A1(n11511), .A2(n16383), .ZN(n8909) );
NOR2_X1 U23904 ( .A1(n11518), .A2(n16383), .ZN(n8761) );
AND2_X1 U23905 ( .A1(n6535), .A2(n1565), .ZN(n6529) );
NOR2_X1 U23906 ( .A1(n11293), .A2(n6536), .ZN(n6535) );
NOR2_X1 U23907 ( .A1(n15797), .A2(n15802), .ZN(n6536) );
NOR2_X1 U23908 ( .A1(n7686), .A2(n7643), .ZN(n7685) );
NOR2_X1 U23909 ( .A1(n7687), .A2(n7688), .ZN(n7686) );
NOR2_X1 U23910 ( .A1(n11147), .A2(n20887), .ZN(n7688) );
NOR2_X1 U23911 ( .A1(n7690), .A2(n7691), .ZN(n7687) );
NOR2_X1 U23912 ( .A1(n9787), .A2(n9788), .ZN(n9786) );
NOR2_X1 U23913 ( .A1(n11145), .A2(n8685), .ZN(n9787) );
NOR2_X1 U23914 ( .A1(n11139), .A2(n8591), .ZN(n9788) );
NOR2_X1 U23915 ( .A1(n8683), .A2(n8684), .ZN(n8682) );
NOR2_X1 U23916 ( .A1(n11309), .A2(n8685), .ZN(n8683) );
NOR2_X1 U23917 ( .A1(n10690), .A2(n16369), .ZN(n8684) );
NOR2_X1 U23918 ( .A1(n9333), .A2(n9334), .ZN(n9332) );
NOR2_X1 U23919 ( .A1(n11148), .A2(n8685), .ZN(n9333) );
NOR2_X1 U23920 ( .A1(n11137), .A2(n8591), .ZN(n9334) );
NOR2_X1 U23921 ( .A1(n9546), .A2(n9547), .ZN(n9545) );
NOR2_X1 U23922 ( .A1(n11483), .A2(n8685), .ZN(n9546) );
NOR2_X1 U23923 ( .A1(n10659), .A2(n8591), .ZN(n9547) );
NOR2_X1 U23924 ( .A1(n8789), .A2(n8790), .ZN(n8788) );
NOR2_X1 U23925 ( .A1(n10695), .A2(n16374), .ZN(n8789) );
NOR2_X1 U23926 ( .A1(n10696), .A2(n16375), .ZN(n8790) );
NOR2_X1 U23927 ( .A1(n8852), .A2(n8853), .ZN(n8851) );
NOR2_X1 U23928 ( .A1(n10677), .A2(n8806), .ZN(n8853) );
NOR2_X1 U23929 ( .A1(n11015), .A2(n16371), .ZN(n8852) );
NAND2_X1 U23930 ( .A1(n4042), .A2(n4043), .ZN(n3427) );
NOR2_X1 U23931 ( .A1(n4057), .A2(n4058), .ZN(n4042) );
NOR2_X1 U23932 ( .A1(n4044), .A2(n4045), .ZN(n4043) );
NOR2_X1 U23933 ( .A1(n10672), .A2(n16355), .ZN(n4058) );
NOR2_X1 U23934 ( .A1(n9066), .A2(n9067), .ZN(n9065) );
NOR2_X1 U23935 ( .A1(n10966), .A2(n16374), .ZN(n9066) );
NOR2_X1 U23936 ( .A1(n10965), .A2(n16375), .ZN(n9067) );
NOR2_X1 U23937 ( .A1(n9107), .A2(n9108), .ZN(n9106) );
NOR2_X1 U23938 ( .A1(n10951), .A2(n16374), .ZN(n9107) );
NOR2_X1 U23939 ( .A1(n10950), .A2(n16375), .ZN(n9108) );
NOR2_X1 U23940 ( .A1(n9148), .A2(n9149), .ZN(n9147) );
NOR2_X1 U23941 ( .A1(n10936), .A2(n16374), .ZN(n9148) );
NOR2_X1 U23942 ( .A1(n10935), .A2(n8567), .ZN(n9149) );
NOR2_X1 U23943 ( .A1(n9189), .A2(n9190), .ZN(n9188) );
NOR2_X1 U23944 ( .A1(n10921), .A2(n16374), .ZN(n9189) );
NOR2_X1 U23945 ( .A1(n10920), .A2(n8567), .ZN(n9190) );
NOR2_X1 U23946 ( .A1(n9230), .A2(n9231), .ZN(n9229) );
NOR2_X1 U23947 ( .A1(n10906), .A2(n16374), .ZN(n9230) );
NOR2_X1 U23948 ( .A1(n10905), .A2(n16375), .ZN(n9231) );
NOR2_X1 U23949 ( .A1(n9271), .A2(n9272), .ZN(n9270) );
NOR2_X1 U23950 ( .A1(n10891), .A2(n16374), .ZN(n9271) );
NOR2_X1 U23951 ( .A1(n10890), .A2(n8567), .ZN(n9272) );
NOR2_X1 U23952 ( .A1(n9369), .A2(n9370), .ZN(n9368) );
AND2_X1 U23953 ( .A1(hart_id_i_20_), .A2(n8581), .ZN(n9370) );
NOR2_X1 U23954 ( .A1(n10885), .A2(n8591), .ZN(n9369) );
NOR2_X1 U23955 ( .A1(n9442), .A2(n9443), .ZN(n9441) );
NOR2_X1 U23956 ( .A1(n10861), .A2(n8572), .ZN(n9442) );
NOR2_X1 U23957 ( .A1(n10860), .A2(n16375), .ZN(n9443) );
NOR2_X1 U23958 ( .A1(n9483), .A2(n9484), .ZN(n9482) );
NOR2_X1 U23959 ( .A1(n10844), .A2(n8572), .ZN(n9483) );
NOR2_X1 U23960 ( .A1(n10843), .A2(n8567), .ZN(n9484) );
NOR2_X1 U23961 ( .A1(n9569), .A2(n9570), .ZN(n9568) );
NOR2_X1 U23962 ( .A1(n10829), .A2(n16374), .ZN(n9569) );
NOR2_X1 U23963 ( .A1(n10828), .A2(n8567), .ZN(n9570) );
NOR2_X1 U23964 ( .A1(n9734), .A2(n9735), .ZN(n9733) );
NOR2_X1 U23965 ( .A1(n11011), .A2(n16371), .ZN(n9734) );
NOR2_X1 U23966 ( .A1(n10768), .A2(n16372), .ZN(n9735) );
NOR2_X1 U23967 ( .A1(n9941), .A2(n9942), .ZN(n9940) );
NOR2_X1 U23968 ( .A1(n11023), .A2(n8590), .ZN(n9942) );
NOR2_X1 U23969 ( .A1(n11008), .A2(n8584), .ZN(n9941) );
NOR2_X1 U23970 ( .A1(n9881), .A2(n9882), .ZN(n9880) );
NOR2_X1 U23971 ( .A1(n11029), .A2(n8590), .ZN(n9882) );
NOR2_X1 U23972 ( .A1(n10661), .A2(n8584), .ZN(n9881) );
NOR2_X1 U23973 ( .A1(n9418), .A2(n9419), .ZN(n9417) );
NOR2_X1 U23974 ( .A1(n11030), .A2(n8590), .ZN(n9419) );
NOR2_X1 U23975 ( .A1(n10644), .A2(n8584), .ZN(n9418) );
NOR2_X1 U23976 ( .A1(n9025), .A2(n9026), .ZN(n9024) );
NOR2_X1 U23977 ( .A1(n11490), .A2(n16374), .ZN(n9025) );
NOR2_X1 U23978 ( .A1(n10637), .A2(n8567), .ZN(n9026) );
NOR2_X1 U23979 ( .A1(n8984), .A2(n8985), .ZN(n8983) );
NOR2_X1 U23980 ( .A1(n10629), .A2(n16374), .ZN(n8984) );
NOR2_X1 U23981 ( .A1(n11491), .A2(n8567), .ZN(n8985) );
NOR2_X1 U23982 ( .A1(n8952), .A2(n8953), .ZN(n8951) );
AND2_X1 U23983 ( .A1(hart_id_i_30_), .A2(n8581), .ZN(n8953) );
NOR2_X1 U23984 ( .A1(n11135), .A2(n16369), .ZN(n8952) );
NAND2_X1 U23985 ( .A1(irq_fast_i_11_), .A2(n16004), .ZN(n7623) );
NAND2_X1 U23986 ( .A1(n9919), .A2(n9920), .ZN(n9900) );
NOR2_X1 U23987 ( .A1(n9928), .A2(n9929), .ZN(n9919) );
NOR2_X1 U23988 ( .A1(n9921), .A2(n9922), .ZN(n9920) );
NOR2_X1 U23989 ( .A1(n11092), .A2(n16362), .ZN(n9929) );
NOR2_X1 U23990 ( .A1(n8582), .A2(n8583), .ZN(n8579) );
NOR2_X1 U23991 ( .A1(n10740), .A2(n8585), .ZN(n8582) );
NOR2_X1 U23992 ( .A1(n10739), .A2(n16372), .ZN(n8583) );
NOR2_X1 U23993 ( .A1(n8629), .A2(n8630), .ZN(n8627) );
NOR2_X1 U23994 ( .A1(n10723), .A2(n16370), .ZN(n8630) );
NOR2_X1 U23995 ( .A1(n10725), .A2(n16372), .ZN(n8629) );
NOR2_X1 U23996 ( .A1(n8718), .A2(n8719), .ZN(n8716) );
NOR2_X1 U23997 ( .A1(n10712), .A2(n8585), .ZN(n8718) );
NOR2_X1 U23998 ( .A1(n10711), .A2(n16372), .ZN(n8719) );
NOR2_X1 U23999 ( .A1(n8791), .A2(n8792), .ZN(n8787) );
NOR2_X1 U24000 ( .A1(n11027), .A2(n16370), .ZN(n8792) );
NOR2_X1 U24001 ( .A1(n10698), .A2(n16372), .ZN(n8791) );
NOR2_X1 U24002 ( .A1(n8854), .A2(n8855), .ZN(n8850) );
NOR2_X1 U24003 ( .A1(n11028), .A2(n16370), .ZN(n8855) );
NOR2_X1 U24004 ( .A1(n10669), .A2(n16372), .ZN(n8854) );
NOR2_X1 U24005 ( .A1(n8902), .A2(n8903), .ZN(n8900) );
NOR2_X1 U24006 ( .A1(n10627), .A2(n8572), .ZN(n8902) );
NOR2_X1 U24007 ( .A1(n11126), .A2(n16375), .ZN(n8903) );
NOR2_X1 U24008 ( .A1(n8745), .A2(n8746), .ZN(n8743) );
NOR2_X1 U24009 ( .A1(n11130), .A2(n8572), .ZN(n8745) );
NOR2_X1 U24010 ( .A1(n11132), .A2(n16375), .ZN(n8746) );
NAND2_X1 U24011 ( .A1(n8705), .A2(n8706), .ZN(n8704) );
NAND2_X1 U24012 ( .A1(n16363), .A2(n16005), .ZN(n8706) );
NOR2_X1 U24013 ( .A1(n8707), .A2(n8708), .ZN(n8705) );
NOR2_X1 U24014 ( .A1(n10709), .A2(n16375), .ZN(n8707) );
NAND2_X1 U24015 ( .A1(irq_fast_i_2_), .A2(n16006), .ZN(n7651) );
NOR2_X1 U24016 ( .A1(n9068), .A2(n9069), .ZN(n9064) );
NOR2_X1 U24017 ( .A1(n10971), .A2(n8590), .ZN(n9069) );
NOR2_X1 U24018 ( .A1(n10975), .A2(n8591), .ZN(n9068) );
NOR2_X1 U24019 ( .A1(n9109), .A2(n9110), .ZN(n9105) );
NOR2_X1 U24020 ( .A1(n10956), .A2(n8590), .ZN(n9110) );
NOR2_X1 U24021 ( .A1(n10960), .A2(n8591), .ZN(n9109) );
NOR2_X1 U24022 ( .A1(n9150), .A2(n9151), .ZN(n9146) );
NOR2_X1 U24023 ( .A1(n10941), .A2(n8590), .ZN(n9151) );
NOR2_X1 U24024 ( .A1(n10945), .A2(n16369), .ZN(n9150) );
NOR2_X1 U24025 ( .A1(n9191), .A2(n9192), .ZN(n9187) );
NOR2_X1 U24026 ( .A1(n10926), .A2(n8590), .ZN(n9192) );
NOR2_X1 U24027 ( .A1(n10930), .A2(n16369), .ZN(n9191) );
NOR2_X1 U24028 ( .A1(n9232), .A2(n9233), .ZN(n9228) );
NOR2_X1 U24029 ( .A1(n10911), .A2(n8590), .ZN(n9233) );
NOR2_X1 U24030 ( .A1(n10915), .A2(n8591), .ZN(n9232) );
NOR2_X1 U24031 ( .A1(n9273), .A2(n9274), .ZN(n9269) );
NOR2_X1 U24032 ( .A1(n10896), .A2(n8590), .ZN(n9274) );
NOR2_X1 U24033 ( .A1(n10900), .A2(n16369), .ZN(n9273) );
NOR2_X1 U24034 ( .A1(n9371), .A2(n9372), .ZN(n9367) );
NOR2_X1 U24035 ( .A1(n10881), .A2(n8590), .ZN(n9372) );
NOR2_X1 U24036 ( .A1(n10878), .A2(n8584), .ZN(n9371) );
NOR2_X1 U24037 ( .A1(n9444), .A2(n9445), .ZN(n9440) );
NOR2_X1 U24038 ( .A1(n10866), .A2(n16370), .ZN(n9445) );
NOR2_X1 U24039 ( .A1(n10870), .A2(n8591), .ZN(n9444) );
NOR2_X1 U24040 ( .A1(n9485), .A2(n9486), .ZN(n9481) );
NOR2_X1 U24041 ( .A1(n10849), .A2(n16370), .ZN(n9486) );
NOR2_X1 U24042 ( .A1(n10853), .A2(n8591), .ZN(n9485) );
NOR2_X1 U24043 ( .A1(n9571), .A2(n9572), .ZN(n9567) );
NOR2_X1 U24044 ( .A1(n10834), .A2(n16370), .ZN(n9572) );
NOR2_X1 U24045 ( .A1(n10838), .A2(n8591), .ZN(n9571) );
NOR2_X1 U24046 ( .A1(n9622), .A2(n9623), .ZN(n9620) );
NOR2_X1 U24047 ( .A1(n10821), .A2(n16371), .ZN(n9622) );
NOR2_X1 U24048 ( .A1(n10816), .A2(n8584), .ZN(n9623) );
NOR2_X1 U24049 ( .A1(n9659), .A2(n9660), .ZN(n9657) );
NOR2_X1 U24050 ( .A1(n10806), .A2(n16371), .ZN(n9659) );
NOR2_X1 U24051 ( .A1(n10802), .A2(n8584), .ZN(n9660) );
NOR2_X1 U24052 ( .A1(n9696), .A2(n9697), .ZN(n9694) );
NOR2_X1 U24053 ( .A1(n10792), .A2(n16371), .ZN(n9696) );
NOR2_X1 U24054 ( .A1(n10787), .A2(n8584), .ZN(n9697) );
NOR2_X1 U24055 ( .A1(n9736), .A2(n9737), .ZN(n9732) );
NOR2_X1 U24056 ( .A1(n10776), .A2(n16370), .ZN(n9737) );
NOR2_X1 U24057 ( .A1(n11138), .A2(n8591), .ZN(n9736) );
NOR2_X1 U24058 ( .A1(n9821), .A2(n9822), .ZN(n9819) );
NOR2_X1 U24059 ( .A1(n10754), .A2(n16371), .ZN(n9821) );
NOR2_X1 U24060 ( .A1(n10753), .A2(n8584), .ZN(n9822) );
NOR2_X1 U24061 ( .A1(n9947), .A2(n9948), .ZN(n9939) );
AND2_X1 U24062 ( .A1(hart_id_i_0_), .A2(n8581), .ZN(n9948) );
NOR2_X1 U24063 ( .A1(n11133), .A2(n8591), .ZN(n9947) );
NOR2_X1 U24064 ( .A1(n9883), .A2(n9884), .ZN(n9879) );
AND2_X1 U24065 ( .A1(hart_id_i_2_), .A2(n8581), .ZN(n9884) );
NOR2_X1 U24066 ( .A1(n11142), .A2(n8591), .ZN(n9883) );
NOR2_X1 U24067 ( .A1(n9420), .A2(n9421), .ZN(n9416) );
AND2_X1 U24068 ( .A1(hart_id_i_1_), .A2(n8581), .ZN(n9421) );
NOR2_X1 U24069 ( .A1(n11143), .A2(n8591), .ZN(n9420) );
NOR2_X1 U24070 ( .A1(n9027), .A2(n9028), .ZN(n9023) );
NOR2_X1 U24071 ( .A1(n10638), .A2(n8590), .ZN(n9028) );
NOR2_X1 U24072 ( .A1(n10642), .A2(n8591), .ZN(n9027) );
NOR2_X1 U24073 ( .A1(n8986), .A2(n8987), .ZN(n8982) );
NOR2_X1 U24074 ( .A1(n11020), .A2(n8590), .ZN(n8987) );
NOR2_X1 U24075 ( .A1(n11136), .A2(n8591), .ZN(n8986) );
NOR2_X1 U24076 ( .A1(n8954), .A2(n8955), .ZN(n8950) );
NOR2_X1 U24077 ( .A1(n11021), .A2(n8590), .ZN(n8955) );
NOR2_X1 U24078 ( .A1(n10615), .A2(n8584), .ZN(n8954) );
NAND2_X1 U24079 ( .A1(n9613), .A2(n9614), .ZN(n9607) );
NOR2_X1 U24080 ( .A1(n15796), .A2(n9615), .ZN(n9614) );
NOR2_X1 U24081 ( .A1(n9616), .A2(n9617), .ZN(n9613) );
NOR2_X1 U24082 ( .A1(n10814), .A2(n8572), .ZN(n9615) );
NAND2_X1 U24083 ( .A1(n9650), .A2(n9651), .ZN(n9644) );
NOR2_X1 U24084 ( .A1(n15796), .A2(n9652), .ZN(n9651) );
NOR2_X1 U24085 ( .A1(n9653), .A2(n9654), .ZN(n9650) );
NOR2_X1 U24086 ( .A1(n10800), .A2(n8572), .ZN(n9652) );
NAND2_X1 U24087 ( .A1(n9687), .A2(n9688), .ZN(n9681) );
NOR2_X1 U24088 ( .A1(n15796), .A2(n9689), .ZN(n9688) );
NOR2_X1 U24089 ( .A1(n9690), .A2(n9691), .ZN(n9687) );
NOR2_X1 U24090 ( .A1(n10785), .A2(n8572), .ZN(n9689) );
NAND2_X1 U24091 ( .A1(n9812), .A2(n9813), .ZN(n9806) );
NOR2_X1 U24092 ( .A1(n15796), .A2(n9814), .ZN(n9813) );
NOR2_X1 U24093 ( .A1(n9815), .A2(n9816), .ZN(n9812) );
NOR2_X1 U24094 ( .A1(n10750), .A2(n8572), .ZN(n9814) );
NAND2_X1 U24095 ( .A1(n1727), .A2(n1728), .ZN(instr_addr_o_5_) );
NAND2_X1 U24096 ( .A1(n15929), .A2(n16007), .ZN(n1728) );
NOR2_X1 U24097 ( .A1(n1730), .A2(n1731), .ZN(n1727) );
NOR2_X1 U24098 ( .A1(n10602), .A2(n1706), .ZN(n1731) );
NOR2_X1 U24099 ( .A1(n9790), .A2(n9791), .ZN(n9785) );
AND2_X1 U24100 ( .A1(hart_id_i_11_), .A2(n8581), .ZN(n9791) );
NOR2_X1 U24101 ( .A1(n11305), .A2(n8688), .ZN(n9790) );
NOR2_X1 U24102 ( .A1(n8686), .A2(n8687), .ZN(n8681) );
AND2_X1 U24103 ( .A1(hart_id_i_7_), .A2(n8581), .ZN(n8687) );
NOR2_X1 U24104 ( .A1(n11476), .A2(n8688), .ZN(n8686) );
NOR2_X1 U24105 ( .A1(n9335), .A2(n9336), .ZN(n9331) );
AND2_X1 U24106 ( .A1(hart_id_i_21_), .A2(n8581), .ZN(n9336) );
NOR2_X1 U24107 ( .A1(n11499), .A2(n8688), .ZN(n9335) );
NOR2_X1 U24108 ( .A1(n9548), .A2(n9549), .ZN(n9544) );
AND2_X1 U24109 ( .A1(hart_id_i_17_), .A2(n8581), .ZN(n9549) );
NOR2_X1 U24110 ( .A1(n10655), .A2(n8688), .ZN(n9548) );
INV_X1 U24111 ( .A(n25148), .ZN(n20088) );
NAND2_X1 U24112 ( .A1(n10347), .A2(n7692), .ZN(n7646) );
NAND2_X1 U24113 ( .A1(irq_fast_i_13_), .A2(n16008), .ZN(n10347) );
NAND2_X1 U24114 ( .A1(irq_fast_i_8_), .A2(n16009), .ZN(n7653) );
NAND2_X1 U24115 ( .A1(n10345), .A2(n7658), .ZN(n7629) );
NAND2_X1 U24116 ( .A1(irq_fast_i_7_), .A2(n16010), .ZN(n10345) );
NAND2_X1 U24117 ( .A1(irq_fast_i_5_), .A2(n16011), .ZN(n7700) );
NAND2_X1 U24118 ( .A1(irq_fast_i_3_), .A2(n16012), .ZN(n7683) );
NAND2_X1 U24119 ( .A1(irq_fast_i_4_), .A2(n16013), .ZN(n7620) );
NAND2_X1 U24120 ( .A1(n11471), .A2(n16439), .ZN(n1706) );
NAND2_X1 U24121 ( .A1(n4034), .A2(n4035), .ZN(n3422) );
NOR2_X1 U24122 ( .A1(n4038), .A2(n4039), .ZN(n4034) );
NOR2_X1 U24123 ( .A1(n4036), .A2(n4037), .ZN(n4035) );
NOR2_X1 U24124 ( .A1(n10703), .A2(n16355), .ZN(n4039) );
NAND2_X1 U24125 ( .A1(n3724), .A2(n3725), .ZN(n3442) );
NOR2_X1 U24126 ( .A1(n3728), .A2(n3729), .ZN(n3724) );
NOR2_X1 U24127 ( .A1(n3726), .A2(n3727), .ZN(n3725) );
NOR2_X1 U24128 ( .A1(n10664), .A2(n16355), .ZN(n3729) );
NAND2_X1 U24129 ( .A1(n4026), .A2(n4027), .ZN(n3417) );
NOR2_X1 U24130 ( .A1(n4030), .A2(n4031), .ZN(n4026) );
NOR2_X1 U24131 ( .A1(n4028), .A2(n4029), .ZN(n4027) );
NOR2_X1 U24132 ( .A1(n11518), .A2(n16355), .ZN(n4031) );
NAND2_X1 U24133 ( .A1(irq_fast_i_12_), .A2(n16014), .ZN(n7692) );
INV_X1 U24134 ( .A(n25140), .ZN(n20140) );
AND2_X1 U24135 ( .A1(n6537), .A2(n11293), .ZN(n6519) );
NOR2_X1 U24136 ( .A1(n20935), .A2(n16462), .ZN(n6537) );
INV_X1 U24137 ( .A(n25170), .ZN(n20030) );
INV_X1 U24138 ( .A(n25169), .ZN(n20086) );
AND2_X1 U24139 ( .A1(n10336), .A2(n7604), .ZN(n7628) );
NAND2_X1 U24140 ( .A1(irq_software_i), .A2(n16015), .ZN(n10336) );
NAND2_X1 U24141 ( .A1(n10152), .A2(n10153), .ZN(n10130) );
NOR2_X1 U24142 ( .A1(n5908), .A2(n10154), .ZN(n10152) );
NAND2_X1 U24143 ( .A1(rf_rdata_b_ecc_i_31_), .A2(n20950), .ZN(n10153) );
NOR2_X1 U24144 ( .A1(n11316), .A2(n5910), .ZN(n10154) );
NAND2_X1 U24145 ( .A1(irq_external_i), .A2(n16016), .ZN(n7604) );
NAND2_X1 U24146 ( .A1(n10918), .A2(n16361), .ZN(n9203) );
NAND2_X1 U24147 ( .A1(n10903), .A2(n16361), .ZN(n9244) );
NAND2_X1 U24148 ( .A1(n10888), .A2(n16361), .ZN(n9285) );
NAND2_X1 U24149 ( .A1(n10858), .A2(n16361), .ZN(n9456) );
NAND2_X1 U24150 ( .A1(n10841), .A2(n16361), .ZN(n9497) );
NAND2_X1 U24151 ( .A1(n10826), .A2(n16361), .ZN(n9583) );
NAND2_X1 U24152 ( .A1(hart_id_i_15_), .A2(n8581), .ZN(n9621) );
NAND2_X1 U24153 ( .A1(hart_id_i_14_), .A2(n8581), .ZN(n9658) );
NAND2_X1 U24154 ( .A1(hart_id_i_13_), .A2(n8581), .ZN(n9695) );
NAND2_X1 U24155 ( .A1(hart_id_i_10_), .A2(n8581), .ZN(n9820) );
NAND2_X1 U24156 ( .A1(hart_id_i_9_), .A2(n8581), .ZN(n8580) );
NAND2_X1 U24157 ( .A1(hart_id_i_6_), .A2(n8581), .ZN(n8717) );
INV_X1 U24158 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_1), .ZN(n20672) );
NAND2_X1 U24159 ( .A1(n5888), .A2(n5889), .ZN(ex_block_i_alu_i_adder_in_b_32) );
NOR2_X1 U24160 ( .A1(n5890), .A2(n5891), .ZN(n5889) );
NOR2_X1 U24161 ( .A1(n5894), .A2(n5895), .ZN(n5888) );
NOR2_X1 U24162 ( .A1(rf_rdata_b_ecc_i_31_), .A2(n20959), .ZN(n5890) );
NAND2_X1 U24163 ( .A1(n11471), .A2(n3018), .ZN(n1708) );
INV_X1 U24164 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_3), .ZN(n20584) );
INV_X1 U24165 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_4), .ZN(n20545) );
INV_X1 U24166 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_2), .ZN(n20638) );
NAND2_X1 U24167 ( .A1(n8845), .A2(n16361), .ZN(n8844) );
OR2_X1 U24168 ( .A1(n8751), .A2(n11151), .ZN(n8845) );
INV_X1 U24169 ( .A(irq_fast_i_7_), .ZN(n20891) );
INV_X1 U24170 ( .A(irq_fast_i_1_), .ZN(n20892) );
INV_X1 U24171 ( .A(irq_timer_i), .ZN(n20882) );
NAND2_X1 U24172 ( .A1(n10963), .A2(n16361), .ZN(n9080) );
NAND2_X1 U24173 ( .A1(n10948), .A2(n16361), .ZN(n9121) );
NAND2_X1 U24174 ( .A1(n10933), .A2(n16361), .ZN(n9162) );
NAND2_X1 U24175 ( .A1(n10694), .A2(n16361), .ZN(n8803) );
NAND2_X1 U24176 ( .A1(n10635), .A2(n16361), .ZN(n9039) );
NAND2_X1 U24177 ( .A1(n10625), .A2(n16361), .ZN(n8998) );
NAND2_X1 U24178 ( .A1(n11510), .A2(n16361), .ZN(n8914) );
NAND2_X1 U24179 ( .A1(n11121), .A2(n16361), .ZN(n8759) );
NAND2_X1 U24180 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U24181 ( .A1(n16471), .A2(n1075), .ZN(n1074) );
NOR2_X1 U24182 ( .A1(n1076), .A2(n1077), .ZN(n1073) );
NOR2_X1 U24183 ( .A1(n11180), .A2(n386), .ZN(n1077) );
NAND2_X1 U24184 ( .A1(n9078), .A2(n9079), .ZN(n9077) );
NOR2_X1 U24185 ( .A1(n9081), .A2(n9082), .ZN(n9078) );
NAND2_X1 U24186 ( .A1(n8758), .A2(n9080), .ZN(n9079) );
NOR2_X1 U24187 ( .A1(n10972), .A2(n8585), .ZN(n9081) );
NAND2_X1 U24188 ( .A1(n9119), .A2(n9120), .ZN(n9118) );
NOR2_X1 U24189 ( .A1(n9122), .A2(n9123), .ZN(n9119) );
NAND2_X1 U24190 ( .A1(n8758), .A2(n9121), .ZN(n9120) );
NOR2_X1 U24191 ( .A1(n10957), .A2(n8585), .ZN(n9122) );
NAND2_X1 U24192 ( .A1(n9160), .A2(n9161), .ZN(n9159) );
NOR2_X1 U24193 ( .A1(n9163), .A2(n9164), .ZN(n9160) );
NAND2_X1 U24194 ( .A1(n8758), .A2(n9162), .ZN(n9161) );
NOR2_X1 U24195 ( .A1(n10942), .A2(n8585), .ZN(n9163) );
NAND2_X1 U24196 ( .A1(n9201), .A2(n9202), .ZN(n9200) );
NOR2_X1 U24197 ( .A1(n9204), .A2(n9205), .ZN(n9201) );
NAND2_X1 U24198 ( .A1(n8758), .A2(n9203), .ZN(n9202) );
NOR2_X1 U24199 ( .A1(n10927), .A2(n8585), .ZN(n9204) );
NAND2_X1 U24200 ( .A1(n9242), .A2(n9243), .ZN(n9241) );
NOR2_X1 U24201 ( .A1(n9245), .A2(n9246), .ZN(n9242) );
NAND2_X1 U24202 ( .A1(n8758), .A2(n9244), .ZN(n9243) );
NOR2_X1 U24203 ( .A1(n10912), .A2(n8585), .ZN(n9245) );
NAND2_X1 U24204 ( .A1(n9283), .A2(n9284), .ZN(n9282) );
NOR2_X1 U24205 ( .A1(n9286), .A2(n9287), .ZN(n9283) );
NAND2_X1 U24206 ( .A1(n8758), .A2(n9285), .ZN(n9284) );
NOR2_X1 U24207 ( .A1(n10897), .A2(n8585), .ZN(n9286) );
NAND2_X1 U24208 ( .A1(n9454), .A2(n9455), .ZN(n9453) );
NOR2_X1 U24209 ( .A1(n9457), .A2(n9458), .ZN(n9454) );
NAND2_X1 U24210 ( .A1(n8758), .A2(n9456), .ZN(n9455) );
NOR2_X1 U24211 ( .A1(n10867), .A2(n16371), .ZN(n9457) );
NAND2_X1 U24212 ( .A1(n9495), .A2(n9496), .ZN(n9494) );
NOR2_X1 U24213 ( .A1(n9498), .A2(n9499), .ZN(n9495) );
NAND2_X1 U24214 ( .A1(n8758), .A2(n9497), .ZN(n9496) );
NOR2_X1 U24215 ( .A1(n10850), .A2(n16371), .ZN(n9498) );
NAND2_X1 U24216 ( .A1(n9581), .A2(n9582), .ZN(n9580) );
NOR2_X1 U24217 ( .A1(n9584), .A2(n9585), .ZN(n9581) );
NAND2_X1 U24218 ( .A1(n8758), .A2(n9583), .ZN(n9582) );
NOR2_X1 U24219 ( .A1(n10835), .A2(n16371), .ZN(n9584) );
NAND2_X1 U24220 ( .A1(n8801), .A2(n8802), .ZN(n8800) );
NOR2_X1 U24221 ( .A1(n8804), .A2(n8805), .ZN(n8801) );
NAND2_X1 U24222 ( .A1(n8758), .A2(n8803), .ZN(n8802) );
NOR2_X1 U24223 ( .A1(n10692), .A2(n8806), .ZN(n8805) );
NAND2_X1 U24224 ( .A1(n9037), .A2(n9038), .ZN(n9036) );
NOR2_X1 U24225 ( .A1(n9040), .A2(n9041), .ZN(n9037) );
NAND2_X1 U24226 ( .A1(n8758), .A2(n9039), .ZN(n9038) );
NOR2_X1 U24227 ( .A1(n10639), .A2(n8585), .ZN(n9040) );
NAND2_X1 U24228 ( .A1(n8996), .A2(n8997), .ZN(n8995) );
NOR2_X1 U24229 ( .A1(n8999), .A2(n9000), .ZN(n8996) );
NAND2_X1 U24230 ( .A1(n8758), .A2(n8998), .ZN(n8997) );
NOR2_X1 U24231 ( .A1(n11494), .A2(n8585), .ZN(n8999) );
NAND2_X1 U24232 ( .A1(n8912), .A2(n8913), .ZN(n8911) );
NOR2_X1 U24233 ( .A1(n8915), .A2(n8916), .ZN(n8912) );
NAND2_X1 U24234 ( .A1(n8758), .A2(n8914), .ZN(n8913) );
NOR2_X1 U24235 ( .A1(n11022), .A2(n16370), .ZN(n8916) );
NAND2_X1 U24236 ( .A1(n8756), .A2(n8757), .ZN(n8755) );
NOR2_X1 U24237 ( .A1(n8760), .A2(n8761), .ZN(n8756) );
NAND2_X1 U24238 ( .A1(n8758), .A2(n8759), .ZN(n8757) );
NOR2_X1 U24239 ( .A1(n11026), .A2(n16370), .ZN(n8760) );
NAND2_X1 U24240 ( .A1(n5896), .A2(n5897), .ZN(n5895) );
NAND2_X1 U24241 ( .A1(n20960), .A2(n11244), .ZN(n5897) );
NAND2_X1 U24242 ( .A1(n20761), .A2(n16409), .ZN(n5896) );
NAND2_X1 U24243 ( .A1(irq_software_i), .A2(n20826), .ZN(n8858) );
NAND2_X1 U24244 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U24245 ( .A1(n78), .A2(n1017), .ZN(n1016) );
NOR2_X1 U24246 ( .A1(n1018), .A2(n1019), .ZN(n1015) );
NOR2_X1 U24247 ( .A1(n11179), .A2(n386), .ZN(n1019) );
NAND2_X1 U24248 ( .A1(n977), .A2(n978), .ZN(n976) );
NAND2_X1 U24249 ( .A1(n78), .A2(n979), .ZN(n978) );
NOR2_X1 U24250 ( .A1(n980), .A2(n981), .ZN(n977) );
NOR2_X1 U24251 ( .A1(n11178), .A2(n386), .ZN(n981) );
NAND2_X1 U24252 ( .A1(n938), .A2(n939), .ZN(n937) );
NAND2_X1 U24253 ( .A1(n16471), .A2(n940), .ZN(n939) );
NOR2_X1 U24254 ( .A1(n941), .A2(n942), .ZN(n938) );
NOR2_X1 U24255 ( .A1(n11177), .A2(n386), .ZN(n942) );
NAND2_X1 U24256 ( .A1(n857), .A2(n858), .ZN(n856) );
NAND2_X1 U24257 ( .A1(n78), .A2(n859), .ZN(n858) );
NOR2_X1 U24258 ( .A1(n860), .A2(n861), .ZN(n857) );
NOR2_X1 U24259 ( .A1(n11176), .A2(n386), .ZN(n861) );
NAND2_X1 U24260 ( .A1(n818), .A2(n819), .ZN(n817) );
NAND2_X1 U24261 ( .A1(n16471), .A2(n820), .ZN(n819) );
NOR2_X1 U24262 ( .A1(n821), .A2(n822), .ZN(n818) );
NOR2_X1 U24263 ( .A1(n11175), .A2(n386), .ZN(n822) );
NAND2_X1 U24264 ( .A1(n780), .A2(n781), .ZN(n779) );
NAND2_X1 U24265 ( .A1(n16471), .A2(n782), .ZN(n781) );
NOR2_X1 U24266 ( .A1(n783), .A2(n784), .ZN(n780) );
NOR2_X1 U24267 ( .A1(n11174), .A2(n386), .ZN(n784) );
NAND2_X1 U24268 ( .A1(n742), .A2(n743), .ZN(n741) );
NAND2_X1 U24269 ( .A1(n16471), .A2(n744), .ZN(n743) );
NOR2_X1 U24270 ( .A1(n745), .A2(n746), .ZN(n742) );
NOR2_X1 U24271 ( .A1(n11173), .A2(n386), .ZN(n746) );
NAND2_X1 U24272 ( .A1(n705), .A2(n706), .ZN(n704) );
NAND2_X1 U24273 ( .A1(n16471), .A2(n707), .ZN(n706) );
NOR2_X1 U24274 ( .A1(n708), .A2(n709), .ZN(n705) );
NOR2_X1 U24275 ( .A1(n11172), .A2(n386), .ZN(n709) );
NAND2_X1 U24276 ( .A1(n667), .A2(n668), .ZN(n666) );
NAND2_X1 U24277 ( .A1(n16471), .A2(n669), .ZN(n668) );
NOR2_X1 U24278 ( .A1(n670), .A2(n671), .ZN(n667) );
NOR2_X1 U24279 ( .A1(n11171), .A2(n386), .ZN(n671) );
NAND2_X1 U24280 ( .A1(n628), .A2(n629), .ZN(n627) );
NAND2_X1 U24281 ( .A1(n16471), .A2(n630), .ZN(n629) );
NOR2_X1 U24282 ( .A1(n631), .A2(n632), .ZN(n628) );
NOR2_X1 U24283 ( .A1(n11170), .A2(n386), .ZN(n632) );
NAND2_X1 U24284 ( .A1(n588), .A2(n589), .ZN(n587) );
NAND2_X1 U24285 ( .A1(n16471), .A2(n590), .ZN(n589) );
NOR2_X1 U24286 ( .A1(n591), .A2(n592), .ZN(n588) );
NOR2_X1 U24287 ( .A1(n11169), .A2(n386), .ZN(n592) );
NAND2_X1 U24288 ( .A1(n548), .A2(n549), .ZN(n547) );
NAND2_X1 U24289 ( .A1(n16471), .A2(n550), .ZN(n549) );
NOR2_X1 U24290 ( .A1(n551), .A2(n552), .ZN(n548) );
NOR2_X1 U24291 ( .A1(n11168), .A2(n386), .ZN(n552) );
NAND2_X1 U24292 ( .A1(n508), .A2(n509), .ZN(n507) );
NAND2_X1 U24293 ( .A1(n16471), .A2(n510), .ZN(n509) );
NOR2_X1 U24294 ( .A1(n511), .A2(n512), .ZN(n508) );
NOR2_X1 U24295 ( .A1(n11167), .A2(n386), .ZN(n512) );
NAND2_X1 U24296 ( .A1(n425), .A2(n426), .ZN(n424) );
NAND2_X1 U24297 ( .A1(n16471), .A2(n427), .ZN(n426) );
NOR2_X1 U24298 ( .A1(n428), .A2(n429), .ZN(n425) );
NOR2_X1 U24299 ( .A1(n11166), .A2(n386), .ZN(n429) );
NAND2_X1 U24300 ( .A1(n9866), .A2(n9362), .ZN(n9865) );
OR2_X1 U24301 ( .A1(n8751), .A2(n11152), .ZN(n9866) );
OR2_X1 U24302 ( .A1(n16270), .A2(n16271), .ZN(n8836) );
NOR2_X1 U24303 ( .A1(n8575), .A2(n11478), .ZN(n16270) );
NOR2_X1 U24304 ( .A1(n16383), .A2(n10672), .ZN(n16271) );
NAND2_X1 U24305 ( .A1(n10342), .A2(n7651), .ZN(n10341) );
NAND2_X1 U24306 ( .A1(irq_fast_i_0_), .A2(n16017), .ZN(n10342) );
INV_X1 U24307 ( .A(n25165), .ZN(n20138) );
NAND2_X1 U24308 ( .A1(n9609), .A2(n9610), .ZN(n9608) );
NAND2_X1 U24309 ( .A1(n16363), .A2(n16018), .ZN(n9610) );
NOR2_X1 U24310 ( .A1(n9611), .A2(n9612), .ZN(n9609) );
NOR2_X1 U24311 ( .A1(n10813), .A2(n8567), .ZN(n9611) );
NAND2_X1 U24312 ( .A1(n9726), .A2(n8621), .ZN(n9718) );
NOR2_X1 U24313 ( .A1(n9728), .A2(n9729), .ZN(n9726) );
NOR2_X1 U24314 ( .A1(n11108), .A2(n16385), .ZN(n9728) );
NOR2_X1 U24315 ( .A1(n11097), .A2(n16362), .ZN(n9729) );
NAND2_X1 U24316 ( .A1(n8620), .A2(n8621), .ZN(n8612) );
NOR2_X1 U24317 ( .A1(n8622), .A2(n8623), .ZN(n8620) );
NOR2_X1 U24318 ( .A1(n10728), .A2(n8102), .ZN(n8622) );
NOR2_X1 U24319 ( .A1(n10727), .A2(n16362), .ZN(n8623) );
NAND2_X1 U24320 ( .A1(n9646), .A2(n9647), .ZN(n9645) );
NAND2_X1 U24321 ( .A1(n16363), .A2(n16019), .ZN(n9647) );
NOR2_X1 U24322 ( .A1(n9648), .A2(n9649), .ZN(n9646) );
NOR2_X1 U24323 ( .A1(n10799), .A2(n8567), .ZN(n9648) );
NAND2_X1 U24324 ( .A1(n9683), .A2(n9684), .ZN(n9682) );
NAND2_X1 U24325 ( .A1(n16363), .A2(n16020), .ZN(n9684) );
NOR2_X1 U24326 ( .A1(n9685), .A2(n9686), .ZN(n9683) );
NOR2_X1 U24327 ( .A1(n10784), .A2(n8567), .ZN(n9685) );
NAND2_X1 U24328 ( .A1(n9808), .A2(n9809), .ZN(n9807) );
NAND2_X1 U24329 ( .A1(n16363), .A2(n16021), .ZN(n9809) );
NOR2_X1 U24330 ( .A1(n9810), .A2(n9811), .ZN(n9808) );
NOR2_X1 U24331 ( .A1(n10749), .A2(n8567), .ZN(n9810) );
NAND2_X1 U24332 ( .A1(n9353), .A2(n9354), .ZN(n9352) );
NOR2_X1 U24333 ( .A1(n9357), .A2(n9358), .ZN(n9353) );
NOR2_X1 U24334 ( .A1(n9355), .A2(n9356), .ZN(n9354) );
NOR2_X1 U24335 ( .A1(n10875), .A2(n8567), .ZN(n9357) );
NAND2_X1 U24336 ( .A1(n8936), .A2(n8937), .ZN(n8935) );
NOR2_X1 U24337 ( .A1(n8940), .A2(n8941), .ZN(n8936) );
NOR2_X1 U24338 ( .A1(n8938), .A2(n8939), .ZN(n8937) );
NOR2_X1 U24339 ( .A1(n11125), .A2(n8567), .ZN(n8940) );
NAND2_X1 U24340 ( .A1(n8568), .A2(n8569), .ZN(n8560) );
NOR2_X1 U24341 ( .A1(n15796), .A2(n8571), .ZN(n8569) );
NOR2_X1 U24342 ( .A1(n8573), .A2(n8574), .ZN(n8568) );
NOR2_X1 U24343 ( .A1(n10735), .A2(n8572), .ZN(n8571) );
NAND2_X1 U24344 ( .A1(n8586), .A2(n8587), .ZN(n8577) );
NOR2_X1 U24345 ( .A1(n8588), .A2(n8589), .ZN(n8587) );
NOR2_X1 U24346 ( .A1(n8592), .A2(n8593), .ZN(n8586) );
NOR2_X1 U24347 ( .A1(n10737), .A2(n16370), .ZN(n8589) );
NAND2_X1 U24348 ( .A1(n8709), .A2(n8710), .ZN(n8703) );
NOR2_X1 U24349 ( .A1(n15796), .A2(n8711), .ZN(n8710) );
NOR2_X1 U24350 ( .A1(n8712), .A2(n8713), .ZN(n8709) );
NOR2_X1 U24351 ( .A1(n10708), .A2(n8572), .ZN(n8711) );
NAND2_X1 U24352 ( .A1(n8720), .A2(n8721), .ZN(n8714) );
NOR2_X1 U24353 ( .A1(n8722), .A2(n8723), .ZN(n8721) );
NOR2_X1 U24354 ( .A1(n8724), .A2(n8725), .ZN(n8720) );
NOR2_X1 U24355 ( .A1(n11025), .A2(n16370), .ZN(n8723) );
NAND2_X1 U24356 ( .A1(n8762), .A2(n8763), .ZN(n8754) );
NOR2_X1 U24357 ( .A1(n8766), .A2(n8767), .ZN(n8762) );
NOR2_X1 U24358 ( .A1(n8764), .A2(n8765), .ZN(n8763) );
AND2_X1 U24359 ( .A1(hart_id_i_5_), .A2(n8581), .ZN(n8766) );
NAND2_X1 U24360 ( .A1(n9083), .A2(n9084), .ZN(n9076) );
NOR2_X1 U24361 ( .A1(n9085), .A2(n9086), .ZN(n9084) );
NOR2_X1 U24362 ( .A1(n9087), .A2(n9088), .ZN(n9083) );
AND2_X1 U24363 ( .A1(hart_id_i_27_), .A2(n8581), .ZN(n9086) );
NAND2_X1 U24364 ( .A1(n9124), .A2(n9125), .ZN(n9117) );
NOR2_X1 U24365 ( .A1(n9126), .A2(n9127), .ZN(n9125) );
NOR2_X1 U24366 ( .A1(n9128), .A2(n9129), .ZN(n9124) );
AND2_X1 U24367 ( .A1(hart_id_i_26_), .A2(n8581), .ZN(n9127) );
NAND2_X1 U24368 ( .A1(n9165), .A2(n9166), .ZN(n9158) );
NOR2_X1 U24369 ( .A1(n9167), .A2(n9168), .ZN(n9166) );
NOR2_X1 U24370 ( .A1(n9169), .A2(n9170), .ZN(n9165) );
AND2_X1 U24371 ( .A1(hart_id_i_25_), .A2(n8581), .ZN(n9168) );
NAND2_X1 U24372 ( .A1(n9206), .A2(n9207), .ZN(n9199) );
NOR2_X1 U24373 ( .A1(n9208), .A2(n9209), .ZN(n9207) );
NOR2_X1 U24374 ( .A1(n9210), .A2(n9211), .ZN(n9206) );
AND2_X1 U24375 ( .A1(hart_id_i_24_), .A2(n8581), .ZN(n9209) );
NAND2_X1 U24376 ( .A1(n9247), .A2(n9248), .ZN(n9240) );
NOR2_X1 U24377 ( .A1(n9249), .A2(n9250), .ZN(n9248) );
NOR2_X1 U24378 ( .A1(n9251), .A2(n9252), .ZN(n9247) );
AND2_X1 U24379 ( .A1(hart_id_i_23_), .A2(n8581), .ZN(n9250) );
NAND2_X1 U24380 ( .A1(n9288), .A2(n9289), .ZN(n9281) );
NOR2_X1 U24381 ( .A1(n9290), .A2(n9291), .ZN(n9289) );
NOR2_X1 U24382 ( .A1(n9292), .A2(n9293), .ZN(n9288) );
AND2_X1 U24383 ( .A1(hart_id_i_22_), .A2(n8581), .ZN(n9291) );
NAND2_X1 U24384 ( .A1(n9459), .A2(n9460), .ZN(n9452) );
NOR2_X1 U24385 ( .A1(n9461), .A2(n9462), .ZN(n9460) );
NOR2_X1 U24386 ( .A1(n9463), .A2(n9464), .ZN(n9459) );
AND2_X1 U24387 ( .A1(hart_id_i_19_), .A2(n8581), .ZN(n9462) );
NAND2_X1 U24388 ( .A1(n9500), .A2(n9501), .ZN(n9493) );
NOR2_X1 U24389 ( .A1(n9502), .A2(n9503), .ZN(n9501) );
NOR2_X1 U24390 ( .A1(n9504), .A2(n9505), .ZN(n9500) );
AND2_X1 U24391 ( .A1(hart_id_i_18_), .A2(n8581), .ZN(n9503) );
NAND2_X1 U24392 ( .A1(n9586), .A2(n9587), .ZN(n9579) );
NOR2_X1 U24393 ( .A1(n9588), .A2(n9589), .ZN(n9587) );
NOR2_X1 U24394 ( .A1(n9590), .A2(n9591), .ZN(n9586) );
AND2_X1 U24395 ( .A1(hart_id_i_16_), .A2(n8581), .ZN(n9589) );
NAND2_X1 U24396 ( .A1(n9042), .A2(n9043), .ZN(n9035) );
NOR2_X1 U24397 ( .A1(n9044), .A2(n9045), .ZN(n9043) );
NOR2_X1 U24398 ( .A1(n9046), .A2(n9047), .ZN(n9042) );
AND2_X1 U24399 ( .A1(hart_id_i_28_), .A2(n8581), .ZN(n9045) );
NAND2_X1 U24400 ( .A1(n9001), .A2(n9002), .ZN(n8994) );
NOR2_X1 U24401 ( .A1(n9003), .A2(n9004), .ZN(n9002) );
NOR2_X1 U24402 ( .A1(n9005), .A2(n9006), .ZN(n9001) );
AND2_X1 U24403 ( .A1(hart_id_i_29_), .A2(n8581), .ZN(n9004) );
NAND2_X1 U24404 ( .A1(n6510), .A2(n6511), .ZN(data_be_o_3_) );
NAND2_X1 U24405 ( .A1(n1564), .A2(n15797), .ZN(n6510) );
NAND2_X1 U24406 ( .A1(n11293), .A2(n6512), .ZN(n6511) );
NAND2_X1 U24407 ( .A1(n6513), .A2(n6514), .ZN(n6512) );
NAND2_X1 U24408 ( .A1(n8917), .A2(n8918), .ZN(n8910) );
NOR2_X1 U24409 ( .A1(n8921), .A2(n8922), .ZN(n8917) );
NOR2_X1 U24410 ( .A1(n8919), .A2(n8920), .ZN(n8918) );
AND2_X1 U24411 ( .A1(hart_id_i_31_), .A2(n8581), .ZN(n8922) );
NAND2_X1 U24412 ( .A1(n9738), .A2(n9739), .ZN(n9730) );
NOR2_X1 U24413 ( .A1(n9742), .A2(n9743), .ZN(n9738) );
NOR2_X1 U24414 ( .A1(n9740), .A2(n9741), .ZN(n9739) );
AND2_X1 U24415 ( .A1(hart_id_i_12_), .A2(n8581), .ZN(n9743) );
NAND2_X1 U24416 ( .A1(n9070), .A2(n9071), .ZN(n9062) );
NOR2_X1 U24417 ( .A1(n9074), .A2(n9075), .ZN(n9070) );
NOR2_X1 U24418 ( .A1(n9072), .A2(n9073), .ZN(n9071) );
NOR2_X1 U24419 ( .A1(n10974), .A2(n16385), .ZN(n9074) );
NAND2_X1 U24420 ( .A1(n9111), .A2(n9112), .ZN(n9103) );
NOR2_X1 U24421 ( .A1(n9115), .A2(n9116), .ZN(n9111) );
NOR2_X1 U24422 ( .A1(n9113), .A2(n9114), .ZN(n9112) );
NOR2_X1 U24423 ( .A1(n10959), .A2(n16385), .ZN(n9115) );
NAND2_X1 U24424 ( .A1(n9152), .A2(n9153), .ZN(n9144) );
NOR2_X1 U24425 ( .A1(n9156), .A2(n9157), .ZN(n9152) );
NOR2_X1 U24426 ( .A1(n9154), .A2(n9155), .ZN(n9153) );
NOR2_X1 U24427 ( .A1(n10944), .A2(n16385), .ZN(n9156) );
NAND2_X1 U24428 ( .A1(n9193), .A2(n9194), .ZN(n9185) );
NOR2_X1 U24429 ( .A1(n9197), .A2(n9198), .ZN(n9193) );
NOR2_X1 U24430 ( .A1(n9195), .A2(n9196), .ZN(n9194) );
NOR2_X1 U24431 ( .A1(n10929), .A2(n16385), .ZN(n9197) );
NAND2_X1 U24432 ( .A1(n9234), .A2(n9235), .ZN(n9226) );
NOR2_X1 U24433 ( .A1(n9238), .A2(n9239), .ZN(n9234) );
NOR2_X1 U24434 ( .A1(n9236), .A2(n9237), .ZN(n9235) );
NOR2_X1 U24435 ( .A1(n10914), .A2(n16385), .ZN(n9238) );
NAND2_X1 U24436 ( .A1(n9275), .A2(n9276), .ZN(n9267) );
NOR2_X1 U24437 ( .A1(n9279), .A2(n9280), .ZN(n9275) );
NOR2_X1 U24438 ( .A1(n9277), .A2(n9278), .ZN(n9276) );
NOR2_X1 U24439 ( .A1(n10899), .A2(n8102), .ZN(n9279) );
NAND2_X1 U24440 ( .A1(n9446), .A2(n9447), .ZN(n9438) );
NOR2_X1 U24441 ( .A1(n9450), .A2(n9451), .ZN(n9446) );
NOR2_X1 U24442 ( .A1(n9448), .A2(n9449), .ZN(n9447) );
NOR2_X1 U24443 ( .A1(n10869), .A2(n16385), .ZN(n9450) );
NAND2_X1 U24444 ( .A1(n9487), .A2(n9488), .ZN(n9479) );
NOR2_X1 U24445 ( .A1(n9491), .A2(n9492), .ZN(n9487) );
NOR2_X1 U24446 ( .A1(n9489), .A2(n9490), .ZN(n9488) );
NOR2_X1 U24447 ( .A1(n10852), .A2(n16385), .ZN(n9491) );
NAND2_X1 U24448 ( .A1(n9573), .A2(n9574), .ZN(n9565) );
NOR2_X1 U24449 ( .A1(n9577), .A2(n9578), .ZN(n9573) );
NOR2_X1 U24450 ( .A1(n9575), .A2(n9576), .ZN(n9574) );
NOR2_X1 U24451 ( .A1(n10837), .A2(n16385), .ZN(n9577) );
NAND2_X1 U24452 ( .A1(n9029), .A2(n9030), .ZN(n9021) );
NOR2_X1 U24453 ( .A1(n9033), .A2(n9034), .ZN(n9029) );
NOR2_X1 U24454 ( .A1(n9031), .A2(n9032), .ZN(n9030) );
NOR2_X1 U24455 ( .A1(n10641), .A2(n16385), .ZN(n9033) );
NAND2_X1 U24456 ( .A1(n8988), .A2(n8989), .ZN(n8980) );
NOR2_X1 U24457 ( .A1(n8992), .A2(n8993), .ZN(n8988) );
NOR2_X1 U24458 ( .A1(n8990), .A2(n8991), .ZN(n8989) );
NOR2_X1 U24459 ( .A1(n11106), .A2(n16385), .ZN(n8992) );
NAND2_X1 U24460 ( .A1(n8904), .A2(n8905), .ZN(n8898) );
NOR2_X1 U24461 ( .A1(n8908), .A2(n8909), .ZN(n8904) );
NOR2_X1 U24462 ( .A1(n8906), .A2(n8907), .ZN(n8905) );
NOR2_X1 U24463 ( .A1(n11104), .A2(n16385), .ZN(n8908) );
NAND2_X1 U24464 ( .A1(n9402), .A2(n9403), .ZN(n9394) );
NOR2_X1 U24465 ( .A1(n9404), .A2(n9405), .ZN(n9403) );
NOR2_X1 U24466 ( .A1(n9406), .A2(n9407), .ZN(n9402) );
NOR2_X1 U24467 ( .A1(n11292), .A2(n8751), .ZN(n9404) );
NAND2_X1 U24468 ( .A1(n8793), .A2(n8794), .ZN(n8785) );
NOR2_X1 U24469 ( .A1(n8797), .A2(n8798), .ZN(n8793) );
NOR2_X1 U24470 ( .A1(n8795), .A2(n8796), .ZN(n8794) );
NOR2_X1 U24471 ( .A1(n10701), .A2(n16385), .ZN(n8797) );
NAND2_X1 U24472 ( .A1(n8747), .A2(n8748), .ZN(n8741) );
NOR2_X1 U24473 ( .A1(n8752), .A2(n8753), .ZN(n8747) );
NOR2_X1 U24474 ( .A1(n8749), .A2(n8750), .ZN(n8748) );
NOR2_X1 U24475 ( .A1(n11110), .A2(n16385), .ZN(n8752) );
NAND2_X1 U24476 ( .A1(n8614), .A2(n8615), .ZN(n8613) );
NOR2_X1 U24477 ( .A1(n8618), .A2(n8619), .ZN(n8614) );
NOR2_X1 U24478 ( .A1(n8616), .A2(n8617), .ZN(n8615) );
NOR2_X1 U24479 ( .A1(n10721), .A2(n8572), .ZN(n8618) );
NAND2_X1 U24480 ( .A1(n8657), .A2(n8658), .ZN(n8656) );
NOR2_X1 U24481 ( .A1(n8661), .A2(n8662), .ZN(n8657) );
NOR2_X1 U24482 ( .A1(n8659), .A2(n8660), .ZN(n8658) );
NOR2_X1 U24483 ( .A1(n10685), .A2(n8572), .ZN(n8661) );
NAND2_X1 U24484 ( .A1(n8673), .A2(n8674), .ZN(n8672) );
NOR2_X1 U24485 ( .A1(n8679), .A2(n8680), .ZN(n8673) );
NOR2_X1 U24486 ( .A1(n8675), .A2(n8676), .ZN(n8674) );
NOR2_X1 U24487 ( .A1(n11024), .A2(n16370), .ZN(n8680) );
NAND2_X1 U24488 ( .A1(n9761), .A2(n9762), .ZN(n9760) );
NOR2_X1 U24489 ( .A1(n9765), .A2(n9766), .ZN(n9761) );
NOR2_X1 U24490 ( .A1(n9763), .A2(n9764), .ZN(n9762) );
NOR2_X1 U24491 ( .A1(n10764), .A2(n8572), .ZN(n9765) );
NAND2_X1 U24492 ( .A1(n9902), .A2(n9903), .ZN(n9901) );
NOR2_X1 U24493 ( .A1(n9911), .A2(n9912), .ZN(n9902) );
NOR2_X1 U24494 ( .A1(n9904), .A2(n9905), .ZN(n9903) );
NOR2_X1 U24495 ( .A1(n11127), .A2(n8572), .ZN(n9911) );
NAND2_X1 U24496 ( .A1(n9856), .A2(n9857), .ZN(n9855) );
NOR2_X1 U24497 ( .A1(n9860), .A2(n9861), .ZN(n9856) );
NOR2_X1 U24498 ( .A1(n9858), .A2(n9859), .ZN(n9857) );
NOR2_X1 U24499 ( .A1(n11129), .A2(n8572), .ZN(n9860) );
NAND2_X1 U24500 ( .A1(n9396), .A2(n9397), .ZN(n9395) );
NOR2_X1 U24501 ( .A1(n9400), .A2(n9401), .ZN(n9396) );
NOR2_X1 U24502 ( .A1(n9398), .A2(n9399), .ZN(n9397) );
NOR2_X1 U24503 ( .A1(n11128), .A2(n16374), .ZN(n9400) );
NAND2_X1 U24504 ( .A1(n9310), .A2(n9311), .ZN(n9309) );
NOR2_X1 U24505 ( .A1(n9314), .A2(n9315), .ZN(n9310) );
NOR2_X1 U24506 ( .A1(n9312), .A2(n9313), .ZN(n9311) );
NOR2_X1 U24507 ( .A1(n11131), .A2(n16374), .ZN(n9314) );
NAND2_X1 U24508 ( .A1(n9522), .A2(n9523), .ZN(n9521) );
NOR2_X1 U24509 ( .A1(n9526), .A2(n9527), .ZN(n9522) );
NOR2_X1 U24510 ( .A1(n9524), .A2(n9525), .ZN(n9523) );
NOR2_X1 U24511 ( .A1(n10653), .A2(n8572), .ZN(n9526) );
NAND2_X1 U24512 ( .A1(n8841), .A2(n8842), .ZN(n8831) );
NOR2_X1 U24513 ( .A1(n8843), .A2(n8844), .ZN(n8842) );
NOR2_X1 U24514 ( .A1(n8846), .A2(n8847), .ZN(n8841) );
NOR2_X1 U24515 ( .A1(n11111), .A2(n16385), .ZN(n8843) );
NAND2_X1 U24516 ( .A1(n8942), .A2(n8943), .ZN(n8934) );
NOR2_X1 U24517 ( .A1(n8944), .A2(n8945), .ZN(n8943) );
NOR2_X1 U24518 ( .A1(n8946), .A2(n8947), .ZN(n8942) );
NOR2_X1 U24519 ( .A1(n11105), .A2(n16385), .ZN(n8944) );
NAND2_X1 U24520 ( .A1(n9359), .A2(n9360), .ZN(n9351) );
NOR2_X1 U24521 ( .A1(n9361), .A2(n8945), .ZN(n9360) );
NOR2_X1 U24522 ( .A1(n9363), .A2(n9364), .ZN(n9359) );
NOR2_X1 U24523 ( .A1(n10884), .A2(n16385), .ZN(n9361) );
NAND2_X1 U24524 ( .A1(n9720), .A2(n9721), .ZN(n9719) );
NOR2_X1 U24525 ( .A1(n9722), .A2(n9723), .ZN(n9721) );
NOR2_X1 U24526 ( .A1(n9724), .A2(n9725), .ZN(n9720) );
NOR2_X1 U24527 ( .A1(n10771), .A2(n16383), .ZN(n9723) );
NAND2_X1 U24528 ( .A1(n9932), .A2(n9933), .ZN(n9931) );
NOR2_X1 U24529 ( .A1(n9936), .A2(n9937), .ZN(n9932) );
NOR2_X1 U24530 ( .A1(n9934), .A2(n9935), .ZN(n9933) );
NOR2_X1 U24531 ( .A1(n10855), .A2(n8806), .ZN(n9937) );
NAND2_X1 U24532 ( .A1(n9776), .A2(n9777), .ZN(n9775) );
NOR2_X1 U24533 ( .A1(n9783), .A2(n9784), .ZN(n9776) );
NOR2_X1 U24534 ( .A1(n9778), .A2(n9779), .ZN(n9777) );
NOR2_X1 U24535 ( .A1(n11018), .A2(n8590), .ZN(n9784) );
NAND2_X1 U24536 ( .A1(n9325), .A2(n9326), .ZN(n9324) );
NOR2_X1 U24537 ( .A1(n9329), .A2(n9330), .ZN(n9325) );
NOR2_X1 U24538 ( .A1(n9327), .A2(n9328), .ZN(n9326) );
NOR2_X1 U24539 ( .A1(n11019), .A2(n8590), .ZN(n9330) );
NAND2_X1 U24540 ( .A1(n9537), .A2(n9538), .ZN(n9536) );
NOR2_X1 U24541 ( .A1(n9542), .A2(n9543), .ZN(n9537) );
NOR2_X1 U24542 ( .A1(n9539), .A2(n9540), .ZN(n9538) );
NOR2_X1 U24543 ( .A1(n10654), .A2(n8590), .ZN(n9543) );
NAND2_X1 U24544 ( .A1(n8631), .A2(n8632), .ZN(n8625) );
NOR2_X1 U24545 ( .A1(n8633), .A2(n8634), .ZN(n8632) );
NOR2_X1 U24546 ( .A1(n8635), .A2(n8636), .ZN(n8631) );
AND2_X1 U24547 ( .A1(hart_id_i_8_), .A2(n8581), .ZN(n8634) );
NAND2_X1 U24548 ( .A1(n8807), .A2(n8808), .ZN(n8799) );
NOR2_X1 U24549 ( .A1(n8809), .A2(n8810), .ZN(n8808) );
NOR2_X1 U24550 ( .A1(n8811), .A2(n8812), .ZN(n8807) );
AND2_X1 U24551 ( .A1(hart_id_i_4_), .A2(n8581), .ZN(n8810) );
NAND2_X1 U24552 ( .A1(n8562), .A2(n8563), .ZN(n8561) );
NAND2_X1 U24553 ( .A1(n16363), .A2(n16022), .ZN(n8563) );
NOR2_X1 U24554 ( .A1(n8565), .A2(n8566), .ZN(n8562) );
NOR2_X1 U24555 ( .A1(n10736), .A2(n16375), .ZN(n8565) );
NAND2_X1 U24556 ( .A1(n9373), .A2(n9374), .ZN(n9365) );
NOR2_X1 U24557 ( .A1(n9377), .A2(n9378), .ZN(n9373) );
NOR2_X1 U24558 ( .A1(n9375), .A2(n9376), .ZN(n9374) );
NOR2_X1 U24559 ( .A1(n10886), .A2(n8685), .ZN(n9377) );
NAND2_X1 U24560 ( .A1(n8956), .A2(n8957), .ZN(n8948) );
NOR2_X1 U24561 ( .A1(n8960), .A2(n8961), .ZN(n8956) );
NOR2_X1 U24562 ( .A1(n8958), .A2(n8959), .ZN(n8957) );
NOR2_X1 U24563 ( .A1(n11146), .A2(n8685), .ZN(n8960) );
NAND2_X1 U24564 ( .A1(n8663), .A2(n8664), .ZN(n8655) );
NOR2_X1 U24565 ( .A1(n8669), .A2(n8670), .ZN(n8663) );
NOR2_X1 U24566 ( .A1(n8665), .A2(n8666), .ZN(n8664) );
NOR2_X1 U24567 ( .A1(n10682), .A2(n16383), .ZN(n8670) );
NAND2_X1 U24568 ( .A1(n9862), .A2(n9863), .ZN(n9854) );
NOR2_X1 U24569 ( .A1(n9869), .A2(n9870), .ZN(n9862) );
NOR2_X1 U24570 ( .A1(n9864), .A2(n9865), .ZN(n9863) );
NOR2_X1 U24571 ( .A1(n11101), .A2(n16362), .ZN(n9870) );
NAND2_X1 U24572 ( .A1(n8833), .A2(n8834), .ZN(n8832) );
NOR2_X1 U24573 ( .A1(n8839), .A2(n8840), .ZN(n8833) );
NOR2_X1 U24574 ( .A1(n8835), .A2(n8836), .ZN(n8834) );
NOR2_X1 U24575 ( .A1(n10674), .A2(n8572), .ZN(n8839) );
INV_X1 U24576 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N37), .ZN(n20639) );
INV_X1 U24577 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N39), .ZN(n20546) );
AND2_X1 U24578 ( .A1(n20826), .A2(irq_external_i), .ZN(n9778) );
AND2_X1 U24579 ( .A1(n20826), .A2(irq_fast_i_5_), .ZN(n9327) );
AND2_X1 U24580 ( .A1(n20826), .A2(irq_fast_i_11_), .ZN(n9088) );
AND2_X1 U24581 ( .A1(n20826), .A2(irq_fast_i_10_), .ZN(n9129) );
AND2_X1 U24582 ( .A1(n20826), .A2(irq_fast_i_9_), .ZN(n9170) );
AND2_X1 U24583 ( .A1(n20826), .A2(irq_fast_i_8_), .ZN(n9211) );
AND2_X1 U24584 ( .A1(n20826), .A2(irq_fast_i_6_), .ZN(n9293) );
AND2_X1 U24585 ( .A1(n20826), .A2(irq_fast_i_4_), .ZN(n9376) );
AND2_X1 U24586 ( .A1(n20826), .A2(irq_fast_i_3_), .ZN(n9464) );
AND2_X1 U24587 ( .A1(n20826), .A2(irq_fast_i_2_), .ZN(n9505) );
AND2_X1 U24588 ( .A1(n20826), .A2(irq_fast_i_0_), .ZN(n9591) );
AND2_X1 U24589 ( .A1(n20826), .A2(irq_fast_i_12_), .ZN(n9047) );
AND2_X1 U24590 ( .A1(n20826), .A2(irq_fast_i_14_), .ZN(n8959) );
INV_X1 U24591 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N38), .ZN(n20585) );
OR2_X1 U24592 ( .A1(n16367), .A2(n10984), .ZN(n8901) );
OR2_X1 U24593 ( .A1(n16368), .A2(n11004), .ZN(n8744) );
OR2_X1 U24594 ( .A1(n8688), .A2(n11477), .ZN(n8862) );
OR2_X1 U24595 ( .A1(n16383), .A2(n10730), .ZN(n8628) );
OR2_X1 U24596 ( .A1(n8856), .A2(n8857), .ZN(n8848) );
NAND2_X1 U24597 ( .A1(n8858), .A2(n8859), .ZN(n8857) );
NAND2_X1 U24598 ( .A1(n8861), .A2(n8862), .ZN(n8856) );
NAND2_X1 U24599 ( .A1(hart_id_i_3_), .A2(n8581), .ZN(n8859) );
NAND2_X1 U24600 ( .A1(n1417), .A2(n1418), .ZN(n1376) );
NAND2_X1 U24601 ( .A1(n1334), .A2(n15886), .ZN(n1417) );
NAND2_X1 U24602 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_0), .A2(n20820), .ZN(n1418) );
NAND2_X1 U24603 ( .A1(n381), .A2(n382), .ZN(n380) );
NAND2_X1 U24604 ( .A1(n16471), .A2(n383), .ZN(n382) );
NOR2_X1 U24605 ( .A1(n384), .A2(n385), .ZN(n381) );
NOR2_X1 U24606 ( .A1(n11216), .A2(n386), .ZN(n385) );
INV_X1 U24607 ( .A(rf_rdata_b_ecc_i_9_), .ZN(n20834) );
INV_X1 U24608 ( .A(rf_rdata_b_ecc_i_8_), .ZN(n20836) );
INV_X1 U24609 ( .A(rf_rdata_b_ecc_i_7_), .ZN(n20840) );
INV_X1 U24610 ( .A(rf_rdata_b_ecc_i_6_), .ZN(n20842) );
INV_X1 U24611 ( .A(rf_rdata_b_ecc_i_5_), .ZN(n20847) );
INV_X1 U24612 ( .A(rf_rdata_b_ecc_i_4_), .ZN(n20854) );
INV_X1 U24613 ( .A(rf_rdata_b_ecc_i_3_), .ZN(n20862) );
INV_X1 U24614 ( .A(rf_rdata_b_ecc_i_2_), .ZN(n20865) );
INV_X1 U24615 ( .A(rf_rdata_b_ecc_i_1_), .ZN(n20870) );
INV_X1 U24616 ( .A(rf_rdata_b_ecc_i_11_), .ZN(n20829) );
INV_X1 U24617 ( .A(rf_rdata_b_ecc_i_10_), .ZN(n20831) );
INV_X1 U24618 ( .A(rf_rdata_b_ecc_i_0_), .ZN(n20872) );
INV_X1 U24619 ( .A(data_rdata_i_7_), .ZN(n20014) );
INV_X1 U24620 ( .A(data_rdata_i_23_), .ZN(n19998) );
INV_X1 U24621 ( .A(data_rdata_i_16_), .ZN(n20005) );
NAND2_X1 U24622 ( .A1(n163), .A2(data_rdata_i_25_), .ZN(n894) );
NAND2_X1 U24623 ( .A1(n163), .A2(data_rdata_i_31_), .ZN(n162) );
NOR2_X1 U24624 ( .A1(n11074), .A2(n16477), .ZN(n879) );
NOR2_X1 U24625 ( .A1(n11075), .A2(n16477), .ZN(n448) );
NOR2_X1 U24626 ( .A1(n11076), .A2(n16477), .ZN(n319) );
NOR2_X1 U24627 ( .A1(n11077), .A2(n44), .ZN(n278) );
NOR2_X1 U24628 ( .A1(n11078), .A2(n44), .ZN(n236) );
NOR2_X1 U24629 ( .A1(n192), .A2(n193), .ZN(n189) );
NOR2_X1 U24630 ( .A1(n11087), .A2(n45), .ZN(n192) );
NOR2_X1 U24631 ( .A1(n11079), .A2(n44), .ZN(n193) );
NOR2_X1 U24632 ( .A1(n144), .A2(n145), .ZN(n141) );
NOR2_X1 U24633 ( .A1(n11088), .A2(n45), .ZN(n144) );
NOR2_X1 U24634 ( .A1(n11080), .A2(n44), .ZN(n145) );
NOR2_X1 U24635 ( .A1(n101), .A2(n102), .ZN(n98) );
NOR2_X1 U24636 ( .A1(n45), .A2(n20021), .ZN(n101) );
NOR2_X1 U24637 ( .A1(n11081), .A2(n44), .ZN(n102) );
NOR2_X1 U24638 ( .A1(n42), .A2(n43), .ZN(n38) );
NOR2_X1 U24639 ( .A1(n45), .A2(n20020), .ZN(n42) );
NOR2_X1 U24640 ( .A1(n11082), .A2(n44), .ZN(n43) );
NOR2_X1 U24641 ( .A1(n648), .A2(n649), .ZN(n646) );
NOR2_X1 U24642 ( .A1(n19996), .A2(n376), .ZN(n648) );
NOR2_X1 U24643 ( .A1(n20012), .A2(n16477), .ZN(n649) );
INV_X1 U24644 ( .A(data_rdata_i_25_), .ZN(n19996) );
INV_X1 U24645 ( .A(data_err_i), .ZN(n20022) );
NOR2_X1 U24646 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U24647 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U24648 ( .A1(n19998), .A2(n72), .ZN(n1111) );
NAND2_X1 U24649 ( .A1(n71), .A2(data_rdata_i_31_), .ZN(n1113) );
NOR2_X1 U24650 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NAND2_X1 U24651 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
NOR2_X1 U24652 ( .A1(n72), .A2(n20003), .ZN(n1321) );
NAND2_X1 U24653 ( .A1(data_rdata_i_26_), .A2(n71), .ZN(n1323) );
NOR2_X1 U24654 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NAND2_X1 U24655 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
NOR2_X1 U24656 ( .A1(n72), .A2(n20002), .ZN(n1267) );
NAND2_X1 U24657 ( .A1(data_rdata_i_27_), .A2(n71), .ZN(n1269) );
NOR2_X1 U24658 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NAND2_X1 U24659 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NOR2_X1 U24660 ( .A1(n72), .A2(n20001), .ZN(n1228) );
NAND2_X1 U24661 ( .A1(data_rdata_i_28_), .A2(n71), .ZN(n1230) );
NOR2_X1 U24662 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U24663 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NOR2_X1 U24664 ( .A1(n72), .A2(n20000), .ZN(n1189) );
NAND2_X1 U24665 ( .A1(data_rdata_i_29_), .A2(n71), .ZN(n1191) );
NOR2_X1 U24666 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND2_X1 U24667 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NOR2_X1 U24668 ( .A1(n72), .A2(n19999), .ZN(n1150) );
NAND2_X1 U24669 ( .A1(data_rdata_i_30_), .A2(n71), .ZN(n1152) );
NOR2_X1 U24670 ( .A1(n459), .A2(n460), .ZN(n458) );
NAND2_X1 U24671 ( .A1(n463), .A2(n464), .ZN(n459) );
NAND2_X1 U24672 ( .A1(n461), .A2(n462), .ZN(n460) );
NAND2_X1 U24673 ( .A1(data_rdata_i_18_), .A2(n21012), .ZN(n464) );
NOR2_X1 U24674 ( .A1(n248), .A2(n249), .ZN(n247) );
NAND2_X1 U24675 ( .A1(n252), .A2(n253), .ZN(n248) );
NAND2_X1 U24676 ( .A1(n250), .A2(n251), .ZN(n249) );
NAND2_X1 U24677 ( .A1(data_rdata_i_21_), .A2(n21012), .ZN(n253) );
NOR2_X1 U24678 ( .A1(n205), .A2(n206), .ZN(n204) );
NAND2_X1 U24679 ( .A1(n209), .A2(n210), .ZN(n205) );
NAND2_X1 U24680 ( .A1(n207), .A2(n208), .ZN(n206) );
NAND2_X1 U24681 ( .A1(data_rdata_i_22_), .A2(n21012), .ZN(n210) );
NOR2_X1 U24682 ( .A1(n159), .A2(n160), .ZN(n158) );
NAND2_X1 U24683 ( .A1(n165), .A2(n166), .ZN(n159) );
NAND2_X1 U24684 ( .A1(n161), .A2(n162), .ZN(n160) );
NAND2_X1 U24685 ( .A1(n21015), .A2(data_rdata_i_15_), .ZN(n165) );
NOR2_X1 U24686 ( .A1(n686), .A2(n687), .ZN(n684) );
NOR2_X1 U24687 ( .A1(n44), .A2(n20013), .ZN(n687) );
NOR2_X1 U24688 ( .A1(n19997), .A2(n376), .ZN(n686) );
INV_X1 U24689 ( .A(data_rdata_i_24_), .ZN(n19997) );
NOR2_X1 U24690 ( .A1(n568), .A2(n569), .ZN(n566) );
NOR2_X1 U24691 ( .A1(n44), .A2(n20010), .ZN(n569) );
NOR2_X1 U24692 ( .A1(n19994), .A2(n376), .ZN(n568) );
INV_X1 U24693 ( .A(data_rdata_i_27_), .ZN(n19994) );
NOR2_X1 U24694 ( .A1(n528), .A2(n529), .ZN(n526) );
NOR2_X1 U24695 ( .A1(n44), .A2(n20009), .ZN(n529) );
NOR2_X1 U24696 ( .A1(n19993), .A2(n376), .ZN(n528) );
INV_X1 U24697 ( .A(data_rdata_i_28_), .ZN(n19993) );
NOR2_X1 U24698 ( .A1(n488), .A2(n489), .ZN(n486) );
NOR2_X1 U24699 ( .A1(n44), .A2(n20008), .ZN(n489) );
NOR2_X1 U24700 ( .A1(n19992), .A2(n376), .ZN(n488) );
INV_X1 U24701 ( .A(data_rdata_i_29_), .ZN(n19992) );
NOR2_X1 U24702 ( .A1(n405), .A2(n406), .ZN(n403) );
NOR2_X1 U24703 ( .A1(n44), .A2(n20007), .ZN(n406) );
NOR2_X1 U24704 ( .A1(n19991), .A2(n376), .ZN(n405) );
INV_X1 U24705 ( .A(data_rdata_i_30_), .ZN(n19991) );
NOR2_X1 U24706 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
NOR2_X1 U24707 ( .A1(n20014), .A2(n45), .ZN(n1095) );
NOR2_X1 U24708 ( .A1(n11088), .A2(n16477), .ZN(n1096) );
NOR2_X1 U24709 ( .A1(n608), .A2(n609), .ZN(n606) );
NOR2_X1 U24710 ( .A1(n44), .A2(n20011), .ZN(n609) );
NOR2_X1 U24711 ( .A1(n376), .A2(n19995), .ZN(n608) );
INV_X1 U24712 ( .A(data_rdata_i_26_), .ZN(n19995) );
NOR2_X1 U24713 ( .A1(n1290), .A2(n1291), .ZN(n1287) );
NOR2_X1 U24714 ( .A1(n45), .A2(n20019), .ZN(n1290) );
NOR2_X1 U24715 ( .A1(n11083), .A2(n16477), .ZN(n1291) );
NOR2_X1 U24716 ( .A1(n1251), .A2(n1252), .ZN(n1248) );
NOR2_X1 U24717 ( .A1(n45), .A2(n20018), .ZN(n1251) );
NOR2_X1 U24718 ( .A1(n11084), .A2(n16477), .ZN(n1252) );
NOR2_X1 U24719 ( .A1(n1212), .A2(n1213), .ZN(n1209) );
NOR2_X1 U24720 ( .A1(n45), .A2(n20017), .ZN(n1212) );
NOR2_X1 U24721 ( .A1(n11085), .A2(n16477), .ZN(n1213) );
NOR2_X1 U24722 ( .A1(n1173), .A2(n1174), .ZN(n1170) );
NOR2_X1 U24723 ( .A1(n45), .A2(n20016), .ZN(n1173) );
NOR2_X1 U24724 ( .A1(n11086), .A2(n16477), .ZN(n1174) );
NOR2_X1 U24725 ( .A1(n1134), .A2(n1135), .ZN(n1131) );
NOR2_X1 U24726 ( .A1(n45), .A2(n20015), .ZN(n1134) );
NOR2_X1 U24727 ( .A1(n11087), .A2(n16477), .ZN(n1135) );
INV_X1 U24728 ( .A(data_rdata_i_21_), .ZN(n20000) );
INV_X1 U24729 ( .A(data_rdata_i_22_), .ZN(n19999) );
INV_X1 U24730 ( .A(data_rdata_i_8_), .ZN(n20013) );
INV_X1 U24731 ( .A(data_rdata_i_15_), .ZN(n20006) );
INV_X1 U24732 ( .A(data_rdata_i_17_), .ZN(n20004) );
INV_X1 U24733 ( .A(data_rdata_i_19_), .ZN(n20002) );
INV_X1 U24734 ( .A(data_rdata_i_20_), .ZN(n20001) );
NAND2_X1 U24735 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U24736 ( .A1(n1051), .A2(n21017), .ZN(n1050) );
NOR2_X1 U24737 ( .A1(n11065), .A2(n1053), .ZN(n1051) );
INV_X1 U24738 ( .A(data_rdata_i_0_), .ZN(n20021) );
INV_X1 U24739 ( .A(data_rdata_i_18_), .ZN(n20003) );
NAND2_X1 U24740 ( .A1(n19966), .A2(data_rdata_i_1_), .ZN(n647) );
NAND2_X1 U24741 ( .A1(data_rdata_i_24_), .A2(n71), .ZN(n120) );
NAND2_X1 U24742 ( .A1(data_rdata_i_25_), .A2(n71), .ZN(n68) );
NAND2_X1 U24743 ( .A1(data_rdata_i_26_), .A2(n163), .ZN(n462) );
NAND2_X1 U24744 ( .A1(data_rdata_i_27_), .A2(n163), .ZN(n334) );
NAND2_X1 U24745 ( .A1(data_rdata_i_28_), .A2(n163), .ZN(n293) );
NAND2_X1 U24746 ( .A1(data_rdata_i_29_), .A2(n163), .ZN(n251) );
NAND2_X1 U24747 ( .A1(data_rdata_i_30_), .A2(n163), .ZN(n208) );
NAND2_X1 U24748 ( .A1(n10306), .A2(n10307), .ZN(n5189) );
NOR2_X1 U24749 ( .A1(n15813), .A2(n15909), .ZN(n10306) );
NOR2_X1 U24750 ( .A1(irq_pending_o), .A2(n10308), .ZN(n10307) );
OR2_X1 U24751 ( .A1(debug_req_i), .A2(irq_nm_i), .ZN(n10308) );
NAND2_X1 U24752 ( .A1(n21014), .A2(data_rdata_i_15_), .ZN(n1056) );
NAND2_X1 U24753 ( .A1(n70), .A2(data_rdata_i_15_), .ZN(n1114) );
INV_X1 U24754 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_0), .ZN(n20681) );
NAND2_X1 U24755 ( .A1(data_rdata_i_0_), .A2(n16346), .ZN(n685) );
NAND2_X1 U24756 ( .A1(data_rdata_i_2_), .A2(n16346), .ZN(n607) );
NAND2_X1 U24757 ( .A1(data_rdata_i_3_), .A2(n16346), .ZN(n567) );
NAND2_X1 U24758 ( .A1(data_rdata_i_4_), .A2(n16346), .ZN(n527) );
NAND2_X1 U24759 ( .A1(data_rdata_i_5_), .A2(n16346), .ZN(n487) );
NAND2_X1 U24760 ( .A1(data_rdata_i_6_), .A2(n16346), .ZN(n404) );
INV_X1 U24761 ( .A(data_rdata_i_9_), .ZN(n20012) );
INV_X1 U24762 ( .A(fetch_enable_i), .ZN(n20895) );
INV_X1 U24763 ( .A(data_rdata_i_31_), .ZN(n19990) );
INV_X1 U24764 ( .A(data_rdata_i_1_), .ZN(n20020) );
INV_X1 U24765 ( .A(data_rdata_i_11_), .ZN(n20010) );
INV_X1 U24766 ( .A(data_rdata_i_12_), .ZN(n20009) );
INV_X1 U24767 ( .A(data_rdata_i_13_), .ZN(n20008) );
INV_X1 U24768 ( .A(data_rdata_i_14_), .ZN(n20007) );
INV_X1 U24769 ( .A(irq_fast_i_13_), .ZN(n20887) );
INV_X1 U24770 ( .A(data_rdata_i_2_), .ZN(n20019) );
INV_X1 U24771 ( .A(data_rdata_i_3_), .ZN(n20018) );
INV_X1 U24772 ( .A(data_rdata_i_4_), .ZN(n20017) );
INV_X1 U24773 ( .A(data_rdata_i_5_), .ZN(n20016) );
INV_X1 U24774 ( .A(data_rdata_i_6_), .ZN(n20015) );
INV_X1 U24775 ( .A(data_rdata_i_10_), .ZN(n20011) );
NAND2_X1 U24776 ( .A1(n4001), .A2(n4002), .ZN(n4000) );
NAND2_X1 U24777 ( .A1(n20925), .A2(n16023), .ZN(n4002) );
NAND2_X1 U24778 ( .A1(boot_addr_i_8_), .A2(n3740), .ZN(n4001) );
NAND2_X1 U24779 ( .A1(n3979), .A2(n3980), .ZN(n3978) );
NAND2_X1 U24780 ( .A1(n20925), .A2(n16024), .ZN(n3980) );
NAND2_X1 U24781 ( .A1(boot_addr_i_10_), .A2(n3740), .ZN(n3979) );
NAND2_X1 U24782 ( .A1(n3956), .A2(n3957), .ZN(n3955) );
NAND2_X1 U24783 ( .A1(n20925), .A2(n16025), .ZN(n3957) );
NAND2_X1 U24784 ( .A1(boot_addr_i_12_), .A2(n3740), .ZN(n3956) );
NAND2_X1 U24785 ( .A1(n3945), .A2(n3946), .ZN(n3944) );
NAND2_X1 U24786 ( .A1(n20925), .A2(n16026), .ZN(n3946) );
NAND2_X1 U24787 ( .A1(boot_addr_i_13_), .A2(n3740), .ZN(n3945) );
NAND2_X1 U24788 ( .A1(n3934), .A2(n3935), .ZN(n3933) );
NAND2_X1 U24789 ( .A1(n20925), .A2(n16027), .ZN(n3935) );
NAND2_X1 U24790 ( .A1(boot_addr_i_14_), .A2(n3740), .ZN(n3934) );
NAND2_X1 U24791 ( .A1(n3923), .A2(n3924), .ZN(n3922) );
NAND2_X1 U24792 ( .A1(n20925), .A2(n16028), .ZN(n3924) );
NAND2_X1 U24793 ( .A1(boot_addr_i_15_), .A2(n3740), .ZN(n3923) );
NAND2_X1 U24794 ( .A1(n3900), .A2(n3901), .ZN(n3899) );
NAND2_X1 U24795 ( .A1(n20925), .A2(n16029), .ZN(n3901) );
NAND2_X1 U24796 ( .A1(boot_addr_i_17_), .A2(n3740), .ZN(n3900) );
NAND2_X1 U24797 ( .A1(n3889), .A2(n3890), .ZN(n3888) );
NAND2_X1 U24798 ( .A1(n20925), .A2(n16030), .ZN(n3890) );
NAND2_X1 U24799 ( .A1(boot_addr_i_18_), .A2(n3740), .ZN(n3889) );
NAND2_X1 U24800 ( .A1(n3878), .A2(n3879), .ZN(n3877) );
NAND2_X1 U24801 ( .A1(n20925), .A2(n16031), .ZN(n3879) );
NAND2_X1 U24802 ( .A1(boot_addr_i_19_), .A2(n16428), .ZN(n3878) );
NAND2_X1 U24803 ( .A1(n3855), .A2(n3856), .ZN(n3854) );
NAND2_X1 U24804 ( .A1(n20925), .A2(n16032), .ZN(n3856) );
NAND2_X1 U24805 ( .A1(boot_addr_i_21_), .A2(n16428), .ZN(n3855) );
NAND2_X1 U24806 ( .A1(n3844), .A2(n3845), .ZN(n3843) );
NAND2_X1 U24807 ( .A1(n20925), .A2(n16033), .ZN(n3845) );
NAND2_X1 U24808 ( .A1(boot_addr_i_22_), .A2(n16428), .ZN(n3844) );
NAND2_X1 U24809 ( .A1(n3833), .A2(n3834), .ZN(n3832) );
NAND2_X1 U24810 ( .A1(n20925), .A2(n16034), .ZN(n3834) );
NAND2_X1 U24811 ( .A1(boot_addr_i_23_), .A2(n16428), .ZN(n3833) );
NAND2_X1 U24812 ( .A1(n3822), .A2(n3823), .ZN(n3821) );
NAND2_X1 U24813 ( .A1(n20925), .A2(n16035), .ZN(n3823) );
NAND2_X1 U24814 ( .A1(boot_addr_i_24_), .A2(n16428), .ZN(n3822) );
NAND2_X1 U24815 ( .A1(n3799), .A2(n3800), .ZN(n3798) );
NAND2_X1 U24816 ( .A1(n20925), .A2(n16036), .ZN(n3800) );
NAND2_X1 U24817 ( .A1(boot_addr_i_26_), .A2(n16428), .ZN(n3799) );
NAND2_X1 U24818 ( .A1(n3760), .A2(n3761), .ZN(n3759) );
NAND2_X1 U24819 ( .A1(n20925), .A2(n16037), .ZN(n3761) );
NAND2_X1 U24820 ( .A1(boot_addr_i_29_), .A2(n16428), .ZN(n3760) );
NAND2_X1 U24821 ( .A1(n3749), .A2(n3750), .ZN(n3748) );
NAND2_X1 U24822 ( .A1(n20925), .A2(n16038), .ZN(n3750) );
NAND2_X1 U24823 ( .A1(boot_addr_i_30_), .A2(n16428), .ZN(n3749) );
NAND2_X1 U24824 ( .A1(n3990), .A2(n3991), .ZN(n3989) );
NAND2_X1 U24825 ( .A1(n20925), .A2(n16039), .ZN(n3991) );
NAND2_X1 U24826 ( .A1(boot_addr_i_9_), .A2(n3740), .ZN(n3990) );
NAND2_X1 U24827 ( .A1(n3736), .A2(n3737), .ZN(n3735) );
NAND2_X1 U24828 ( .A1(n20925), .A2(n16040), .ZN(n3737) );
NAND2_X1 U24829 ( .A1(boot_addr_i_31_), .A2(n3740), .ZN(n3736) );
INV_X1 U24830 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N35), .ZN(n20682) );
NAND2_X1 U24831 ( .A1(n21015), .A2(data_rdata_i_9_), .ZN(n895) );
NAND2_X1 U24832 ( .A1(n21012), .A2(data_rdata_i_17_), .ZN(n896) );
NAND2_X1 U24833 ( .A1(n21012), .A2(data_rdata_i_23_), .ZN(n166) );
INV_X1 U24834 ( .A(data_rvalid_i), .ZN(n19989) );
NAND2_X1 U24835 ( .A1(n875), .A2(n876), .ZN(n874) );
NOR2_X1 U24836 ( .A1(n878), .A2(n879), .ZN(n875) );
NAND2_X1 U24837 ( .A1(n19966), .A2(n16080), .ZN(n876) );
NOR2_X1 U24838 ( .A1(n11082), .A2(n45), .ZN(n878) );
NAND2_X1 U24839 ( .A1(n444), .A2(n445), .ZN(n443) );
NOR2_X1 U24840 ( .A1(n447), .A2(n448), .ZN(n444) );
NAND2_X1 U24841 ( .A1(n19966), .A2(n16079), .ZN(n445) );
NOR2_X1 U24842 ( .A1(n11083), .A2(n45), .ZN(n447) );
NAND2_X1 U24843 ( .A1(data_rdata_i_8_), .A2(n70), .ZN(n121) );
NAND2_X1 U24844 ( .A1(data_rdata_i_9_), .A2(n70), .ZN(n69) );
NAND2_X1 U24845 ( .A1(data_rdata_i_10_), .A2(n70), .ZN(n1324) );
NAND2_X1 U24846 ( .A1(data_rdata_i_11_), .A2(n70), .ZN(n1270) );
NAND2_X1 U24847 ( .A1(data_rdata_i_12_), .A2(n70), .ZN(n1231) );
NAND2_X1 U24848 ( .A1(data_rdata_i_13_), .A2(n70), .ZN(n1192) );
NAND2_X1 U24849 ( .A1(data_rdata_i_14_), .A2(n70), .ZN(n1153) );
NAND2_X1 U24850 ( .A1(n315), .A2(n316), .ZN(n314) );
NAND2_X1 U24851 ( .A1(n16346), .A2(n16078), .ZN(n316) );
NOR2_X1 U24852 ( .A1(n318), .A2(n319), .ZN(n315) );
NOR2_X1 U24853 ( .A1(n11084), .A2(n45), .ZN(n318) );
NAND2_X1 U24854 ( .A1(n274), .A2(n275), .ZN(n273) );
NAND2_X1 U24855 ( .A1(n16346), .A2(n16077), .ZN(n275) );
NOR2_X1 U24856 ( .A1(n277), .A2(n278), .ZN(n274) );
NOR2_X1 U24857 ( .A1(n11085), .A2(n45), .ZN(n277) );
NAND2_X1 U24858 ( .A1(n232), .A2(n233), .ZN(n231) );
NAND2_X1 U24859 ( .A1(n16346), .A2(n16076), .ZN(n233) );
NOR2_X1 U24860 ( .A1(n235), .A2(n236), .ZN(n232) );
NOR2_X1 U24861 ( .A1(n11086), .A2(n45), .ZN(n235) );
NAND2_X1 U24862 ( .A1(data_rdata_i_1_), .A2(n21014), .ZN(n893) );
NAND2_X1 U24863 ( .A1(data_rdata_i_2_), .A2(n21014), .ZN(n461) );
NAND2_X1 U24864 ( .A1(data_rdata_i_3_), .A2(n21014), .ZN(n333) );
NAND2_X1 U24865 ( .A1(data_rdata_i_4_), .A2(n21014), .ZN(n292) );
NAND2_X1 U24866 ( .A1(data_rdata_i_5_), .A2(n21014), .ZN(n250) );
NAND2_X1 U24867 ( .A1(data_rdata_i_6_), .A2(n21014), .ZN(n207) );
NAND2_X1 U24868 ( .A1(data_rdata_i_7_), .A2(n21014), .ZN(n161) );
NAND2_X1 U24869 ( .A1(boot_addr_i_11_), .A2(n3740), .ZN(n3972) );
NAND2_X1 U24870 ( .A1(boot_addr_i_16_), .A2(n3740), .ZN(n3916) );
NAND2_X1 U24871 ( .A1(boot_addr_i_20_), .A2(n16428), .ZN(n3871) );
NAND2_X1 U24872 ( .A1(boot_addr_i_25_), .A2(n16428), .ZN(n3815) );
NAND2_X1 U24873 ( .A1(boot_addr_i_27_), .A2(n16428), .ZN(n3792) );
NAND2_X1 U24874 ( .A1(boot_addr_i_28_), .A2(n16428), .ZN(n3780) );
NAND2_X1 U24875 ( .A1(data_rdata_i_19_), .A2(n21012), .ZN(n336) );
NAND2_X1 U24876 ( .A1(data_rdata_i_20_), .A2(n21012), .ZN(n295) );
AND2_X1 U24877 ( .A1(data_rdata_i_24_), .A2(n163), .ZN(n1362) );
NAND2_X1 U24878 ( .A1(data_rdata_i_10_), .A2(n21015), .ZN(n463) );
NAND2_X1 U24879 ( .A1(data_rdata_i_11_), .A2(n21015), .ZN(n335) );
NAND2_X1 U24880 ( .A1(data_rdata_i_12_), .A2(n21015), .ZN(n294) );
NAND2_X1 U24881 ( .A1(data_rdata_i_13_), .A2(n21015), .ZN(n252) );
NAND2_X1 U24882 ( .A1(data_rdata_i_14_), .A2(n21015), .ZN(n209) );
NAND2_X1 U24883 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
OR2_X1 U24884 ( .A1(n16477), .A2(n11073), .ZN(n1348) );
NAND2_X1 U24885 ( .A1(n19966), .A2(n16057), .ZN(n1347) );
NOR2_X1 U24886 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U24887 ( .A1(n1059), .A2(n1060), .ZN(n1054) );
NAND2_X1 U24888 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U24889 ( .A1(data_rdata_i_31_), .A2(n21013), .ZN(n1060) );
OR2_X1 U24890 ( .A1(n45), .A2(n11081), .ZN(n1352) );
NAND2_X1 U24891 ( .A1(n1298), .A2(n1299), .ZN(n1049) );
NOR2_X1 U24892 ( .A1(n11064), .A2(n11065), .ZN(n1298) );
NAND2_X1 U24893 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
NOR2_X1 U24894 ( .A1(n1306), .A2(n1307), .ZN(n1300) );
NAND2_X1 U24895 ( .A1(n21016), .A2(data_rdata_i_23_), .ZN(n1059) );
NAND2_X1 U24896 ( .A1(n7024), .A2(n7019), .ZN(n6712) );
NOR2_X1 U24897 ( .A1(n11345), .A2(n7025), .ZN(n7024) );
NOR2_X1 U24898 ( .A1(n11153), .A2(n5712), .ZN(n5710) );
AND2_X1 U24899 ( .A1(n5273), .A2(n5532), .ZN(n5712) );
NOR2_X1 U24900 ( .A1(instr_rvalid_i), .A2(n15920), .ZN(n3721) );
NOR2_X1 U24901 ( .A1(n11519), .A2(n11520), .ZN(n5238) );
NOR2_X1 U24902 ( .A1(n2848), .A2(n2849), .ZN(n2844) );
NOR2_X1 U24903 ( .A1(n2846), .A2(n2847), .ZN(n2845) );
NOR2_X1 U24904 ( .A1(n11367), .A2(n2169), .ZN(n2848) );
NOR2_X1 U24905 ( .A1(n11519), .A2(n5221), .ZN(n10448) );
NAND2_X1 U24906 ( .A1(n3575), .A2(n3576), .ZN(n3290) );
NOR2_X1 U24907 ( .A1(n3584), .A2(n3585), .ZN(n3575) );
NOR2_X1 U24908 ( .A1(n3577), .A2(n3578), .ZN(n3576) );
NOR2_X1 U24909 ( .A1(n11460), .A2(n16450), .ZN(n3585) );
NAND2_X1 U24910 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_1), .ZN(n22097) );
NAND2_X1 U24911 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_1), .A2(n11254), .ZN(n22094) );
NAND2_X1 U24912 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_2), .A2(n11255), .ZN(n22095) );
NOR2_X1 U24913 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_0), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_N218), .ZN(n5010) );
NAND2_X1 U24914 ( .A1(n11459), .A2(crash_dump_o_65_), .ZN(n2166) );
AND2_X1 U24915 ( .A1(n6187), .A2(n6188), .ZN(n6077) );
NAND2_X1 U24916 ( .A1(n20953), .A2(n6190), .ZN(n6188) );
NOR2_X1 U24917 ( .A1(n11316), .A2(n16356), .ZN(n6187) );
NAND2_X1 U24918 ( .A1(n22105), .A2(n22104), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_N219) );
NAND2_X1 U24919 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_2), .A2(n22103), .ZN(n22104) );
NOR2_X1 U24920 ( .A1(n6540), .A2(n11313), .ZN(n1590) );
NOR2_X1 U24921 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fifo_i_add_146_B_1_), .A2(n11485), .ZN(n21446) );
NAND2_X1 U24922 ( .A1(n2879), .A2(n2880), .ZN(n2440) );
NOR2_X1 U24923 ( .A1(n2884), .A2(n2885), .ZN(n2879) );
NOR2_X1 U24924 ( .A1(n2881), .A2(n2882), .ZN(n2880) );
NOR2_X1 U24925 ( .A1(n11369), .A2(n16448), .ZN(n2884) );
NOR2_X1 U24926 ( .A1(n11341), .A2(n11343), .ZN(n10230) );
NAND2_X1 U24927 ( .A1(n11468), .A2(n3019), .ZN(n3042) );
NAND2_X1 U24928 ( .A1(n2887), .A2(n2888), .ZN(n2035) );
NOR2_X1 U24929 ( .A1(n2892), .A2(n2893), .ZN(n2887) );
NOR2_X1 U24930 ( .A1(n2889), .A2(n2890), .ZN(n2888) );
NOR2_X1 U24931 ( .A1(n11373), .A2(n16448), .ZN(n2892) );
NAND2_X1 U24932 ( .A1(n11517), .A2(n10464), .ZN(n4056) );
NAND2_X1 U24933 ( .A1(n2838), .A2(n2839), .ZN(n2275) );
NOR2_X1 U24934 ( .A1(n2842), .A2(n2843), .ZN(n2838) );
NOR2_X1 U24935 ( .A1(n2840), .A2(n2841), .ZN(n2839) );
NOR2_X1 U24936 ( .A1(n11461), .A2(n16448), .ZN(n2842) );
NAND2_X1 U24937 ( .A1(n1549), .A2(n1598), .ZN(n1507) );
NAND2_X1 U24938 ( .A1(n1599), .A2(n1571), .ZN(n1598) );
NAND2_X1 U24939 ( .A1(n1579), .A2(n1600), .ZN(n1599) );
NAND2_X1 U24940 ( .A1(n11298), .A2(n1601), .ZN(n1600) );
NAND2_X1 U24941 ( .A1(n2852), .A2(n2853), .ZN(n2103) );
NOR2_X1 U24942 ( .A1(n2856), .A2(n2857), .ZN(n2852) );
NOR2_X1 U24943 ( .A1(n2854), .A2(n2855), .ZN(n2853) );
NOR2_X1 U24944 ( .A1(n11365), .A2(n16448), .ZN(n2856) );
NOR2_X1 U24945 ( .A1(n1447), .A2(n1448), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fifo_i_add_146_B_1_) );
NOR2_X1 U24946 ( .A1(n1449), .A2(n11485), .ZN(n1448) );
NOR2_X1 U24947 ( .A1(n20111), .A2(n16197), .ZN(n5541) );
NOR2_X1 U24948 ( .A1(n10253), .A2(n11339), .ZN(n10099) );
NAND2_X1 U24949 ( .A1(n10298), .A2(n20965), .ZN(n10185) );
NOR2_X1 U24950 ( .A1(n11326), .A2(n15799), .ZN(n10298) );
NAND2_X1 U24951 ( .A1(n2806), .A2(n2807), .ZN(n2136) );
NOR2_X1 U24952 ( .A1(n2811), .A2(n2812), .ZN(n2806) );
NOR2_X1 U24953 ( .A1(n2808), .A2(n2809), .ZN(n2807) );
NOR2_X1 U24954 ( .A1(n11355), .A2(n16448), .ZN(n2811) );
NOR2_X1 U24955 ( .A1(n11290), .A2(n11289), .ZN(n4426) );
NAND2_X1 U24956 ( .A1(n11297), .A2(n19965), .ZN(n1549) );
NAND2_X1 U24957 ( .A1(n2798), .A2(n2799), .ZN(n2018) );
NOR2_X1 U24958 ( .A1(n2803), .A2(n2804), .ZN(n2798) );
NOR2_X1 U24959 ( .A1(n2800), .A2(n2801), .ZN(n2799) );
NOR2_X1 U24960 ( .A1(n11357), .A2(n2169), .ZN(n2803) );
NAND2_X1 U24961 ( .A1(n11319), .A2(n15893), .ZN(n10182) );
NAND2_X1 U24962 ( .A1(n7721), .A2(n11498), .ZN(n7023) );
AND2_X1 U24963 ( .A1(n7722), .A2(n7716), .ZN(n7721) );
NAND2_X1 U24964 ( .A1(n11501), .A2(n15804), .ZN(n1440) );
NAND2_X1 U24965 ( .A1(n2864), .A2(n2865), .ZN(n2727) );
NOR2_X1 U24966 ( .A1(n2868), .A2(n2869), .ZN(n2864) );
NOR2_X1 U24967 ( .A1(n2866), .A2(n2867), .ZN(n2865) );
NOR2_X1 U24968 ( .A1(n11391), .A2(n2169), .ZN(n2868) );
NAND2_X1 U24969 ( .A1(n22107), .A2(n22106), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_N220) );
NAND2_X1 U24970 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_3), .A2(n22105), .ZN(n22106) );
NAND2_X1 U24971 ( .A1(n2789), .A2(n2790), .ZN(n2203) );
NOR2_X1 U24972 ( .A1(n2794), .A2(n2795), .ZN(n2789) );
NOR2_X1 U24973 ( .A1(n2791), .A2(n2792), .ZN(n2790) );
NOR2_X1 U24974 ( .A1(n11351), .A2(n16448), .ZN(n2794) );
NAND2_X1 U24975 ( .A1(n22103), .A2(n22102), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_N218) );
NAND2_X1 U24976 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_1), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_0), .ZN(n22102) );
NAND2_X1 U24977 ( .A1(n11300), .A2(n15922), .ZN(n4958) );
NOR2_X1 U24978 ( .A1(n2525), .A2(n2526), .ZN(n2519) );
AND2_X1 U24979 ( .A1(n2530), .A2(n2531), .ZN(n2525) );
NAND2_X1 U24980 ( .A1(n2527), .A2(n2528), .ZN(n2526) );
NAND2_X1 U24981 ( .A1(n11405), .A2(n15803), .ZN(n2531) );
NAND2_X1 U24982 ( .A1(n3601), .A2(n3594), .ZN(n3050) );
NOR2_X1 U24983 ( .A1(n3603), .A2(n3604), .ZN(n3601) );
NOR2_X1 U24984 ( .A1(n11460), .A2(n3605), .ZN(n3604) );
NOR2_X1 U24985 ( .A1(n19960), .A2(n3606), .ZN(n3603) );
NOR2_X1 U24986 ( .A1(n1554), .A2(data_rvalid_i), .ZN(n1528) );
NOR2_X1 U24987 ( .A1(n1501), .A2(data_gnt_i), .ZN(n1548) );
NAND2_X1 U24988 ( .A1(n10467), .A2(n10468), .ZN(n5221) );
NOR2_X1 U24989 ( .A1(n15798), .A2(n15819), .ZN(n10467) );
NOR2_X1 U24990 ( .A1(n11516), .A2(n11517), .ZN(n10468) );
NAND2_X1 U24991 ( .A1(n11502), .A2(n15895), .ZN(n1442) );
NAND2_X1 U24992 ( .A1(n6302), .A2(n11290), .ZN(n4941) );
NOR2_X1 U24993 ( .A1(n11289), .A2(n15888), .ZN(n6302) );
NOR2_X1 U24994 ( .A1(n11475), .A2(n3028), .ZN(n3025) );
AND2_X1 U24995 ( .A1(n21491), .A2(crash_dump_o_67_), .ZN(n21486) );
NOR2_X1 U24996 ( .A1(n11313), .A2(n11320), .ZN(n10290) );
NOR2_X1 U24997 ( .A1(n11519), .A2(n11301), .ZN(n5133) );
INV_X1 U24998 ( .A(instr_rdata_i_1_), .ZN(n19960) );
NAND2_X1 U24999 ( .A1(n5375), .A2(n5376), .ZN(n4435) );
NAND2_X1 U25000 ( .A1(n5377), .A2(n15891), .ZN(n5376) );
NAND2_X1 U25001 ( .A1(n11244), .A2(n20112), .ZN(n5375) );
NAND2_X1 U25002 ( .A1(data_addr_o_31_), .A2(n16041), .ZN(n5377) );
NOR2_X1 U25003 ( .A1(n2746), .A2(n3602), .ZN(n3594) );
NOR2_X1 U25004 ( .A1(n11460), .A2(n11390), .ZN(n3602) );
NOR2_X1 U25005 ( .A1(n11253), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_4), .ZN(n22086) );
NAND2_X1 U25006 ( .A1(n20991), .A2(n8142), .ZN(n7722) );
NAND2_X1 U25007 ( .A1(n15800), .A2(n8143), .ZN(n8142) );
NAND2_X1 U25008 ( .A1(n11498), .A2(n5196), .ZN(n8143) );
NOR2_X1 U25009 ( .A1(n15911), .A2(n1372), .ZN(n1365) );
NAND2_X1 U25010 ( .A1(n11294), .A2(n11297), .ZN(n1372) );
NOR2_X1 U25011 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_4), .ZN(n22088) );
NAND2_X1 U25012 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_0), .A2(n22086), .ZN(n22101) );
NAND2_X1 U25013 ( .A1(n22088), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_0), .ZN(n22098) );
NAND2_X1 U25014 ( .A1(n22087), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_0), .ZN(n22090) );
NAND2_X1 U25015 ( .A1(n22091), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_0), .ZN(n22093) );
NAND2_X1 U25016 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N218), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_0), .ZN(n4996) );
NAND2_X1 U25017 ( .A1(n11062), .A2(n11091), .ZN(n1040) );
NAND2_X1 U25018 ( .A1(n11091), .A2(n15923), .ZN(n1305) );
NAND2_X1 U25019 ( .A1(n10537), .A2(n11295), .ZN(n1571) );
NOR2_X1 U25020 ( .A1(n11296), .A2(n11298), .ZN(n10537) );
NAND2_X1 U25021 ( .A1(n8422), .A2(n20993), .ZN(n5116) );
NOR2_X1 U25022 ( .A1(n19988), .A2(n8424), .ZN(n8422) );
NOR2_X1 U25023 ( .A1(n16131), .A2(n1698), .ZN(n8424) );
NAND2_X1 U25024 ( .A1(n10367), .A2(n11313), .ZN(n10374) );
NAND2_X1 U25025 ( .A1(n10295), .A2(n10296), .ZN(n4939) );
NOR2_X1 U25026 ( .A1(n11328), .A2(n15914), .ZN(n10296) );
NOR2_X1 U25027 ( .A1(n10185), .A2(n5583), .ZN(n10295) );
NAND2_X1 U25028 ( .A1(n11289), .A2(n11291), .ZN(n5556) );
NAND2_X1 U25029 ( .A1(n2817), .A2(n2818), .ZN(n2051) );
NOR2_X1 U25030 ( .A1(n2821), .A2(n2822), .ZN(n2817) );
NOR2_X1 U25031 ( .A1(n2819), .A2(n2820), .ZN(n2818) );
NOR2_X1 U25032 ( .A1(n11359), .A2(n2169), .ZN(n2821) );
NAND2_X1 U25033 ( .A1(n11297), .A2(n19989), .ZN(n1580) );
NOR2_X1 U25034 ( .A1(n11492), .A2(n6793), .ZN(n6820) );
NOR2_X1 U25035 ( .A1(n11051), .A2(n6793), .ZN(n6892) );
NOR2_X1 U25036 ( .A1(n11057), .A2(n6793), .ZN(n6838) );
NOR2_X1 U25037 ( .A1(n11056), .A2(n6793), .ZN(n6847) );
NOR2_X1 U25038 ( .A1(n11055), .A2(n6793), .ZN(n6856) );
NOR2_X1 U25039 ( .A1(n11054), .A2(n6793), .ZN(n6865) );
NOR2_X1 U25040 ( .A1(n11053), .A2(n6793), .ZN(n6874) );
NOR2_X1 U25041 ( .A1(n11052), .A2(n6793), .ZN(n6883) );
NOR2_X1 U25042 ( .A1(n11050), .A2(n6793), .ZN(n6901) );
NOR2_X1 U25043 ( .A1(n11049), .A2(n6793), .ZN(n6921) );
NOR2_X1 U25044 ( .A1(n11048), .A2(n6793), .ZN(n6930) );
NOR2_X1 U25045 ( .A1(n11046), .A2(n6793), .ZN(n6948) );
NOR2_X1 U25046 ( .A1(n11047), .A2(n6793), .ZN(n6939) );
NOR2_X1 U25047 ( .A1(n11058), .A2(n6793), .ZN(n6829) );
NOR2_X1 U25048 ( .A1(n11059), .A2(n6793), .ZN(n6799) );
NOR2_X1 U25049 ( .A1(n11060), .A2(n6793), .ZN(n6787) );
NOR2_X1 U25050 ( .A1(n11493), .A2(n6796), .ZN(n6825) );
NOR2_X1 U25051 ( .A1(n11331), .A2(n6796), .ZN(n6897) );
NOR2_X1 U25052 ( .A1(n11336), .A2(n6796), .ZN(n6843) );
NOR2_X1 U25053 ( .A1(n11334), .A2(n6796), .ZN(n6852) );
NOR2_X1 U25054 ( .A1(n11325), .A2(n6796), .ZN(n6861) );
NOR2_X1 U25055 ( .A1(n11311), .A2(n6796), .ZN(n6870) );
NOR2_X1 U25056 ( .A1(n11332), .A2(n6796), .ZN(n6879) );
NOR2_X1 U25057 ( .A1(n11323), .A2(n6796), .ZN(n6888) );
NOR2_X1 U25058 ( .A1(n11330), .A2(n6796), .ZN(n6906) );
NOR2_X1 U25059 ( .A1(n11338), .A2(n6796), .ZN(n6834) );
NOR2_X1 U25060 ( .A1(n11340), .A2(n6796), .ZN(n6804) );
NOR2_X1 U25061 ( .A1(n11316), .A2(n6796), .ZN(n6794) );
NAND2_X1 U25062 ( .A1(n2858), .A2(n2859), .ZN(n2432) );
NAND2_X1 U25063 ( .A1(n16449), .A2(n15821), .ZN(n2859) );
NOR2_X1 U25064 ( .A1(n2861), .A2(n2862), .ZN(n2858) );
NOR2_X1 U25065 ( .A1(n11485), .A2(n19943), .ZN(n2861) );
NAND2_X1 U25066 ( .A1(n2776), .A2(n2777), .ZN(n2426) );
NOR2_X1 U25067 ( .A1(n2780), .A2(n2781), .ZN(n2776) );
NOR2_X1 U25068 ( .A1(n2778), .A2(n2779), .ZN(n2777) );
NOR2_X1 U25069 ( .A1(n11353), .A2(n16448), .ZN(n2780) );
NOR2_X1 U25070 ( .A1(n11389), .A2(n2756), .ZN(n2889) );
NOR2_X1 U25071 ( .A1(n11388), .A2(n2756), .ZN(n2873) );
NOR2_X1 U25072 ( .A1(n11462), .A2(n2756), .ZN(n2840) );
NOR2_X1 U25073 ( .A1(n11387), .A2(n2756), .ZN(n2881) );
NOR2_X1 U25074 ( .A1(n11381), .A2(n2756), .ZN(n2800) );
NOR2_X1 U25075 ( .A1(n11386), .A2(n2756), .ZN(n2846) );
NOR2_X1 U25076 ( .A1(n11383), .A2(n2756), .ZN(n2832) );
NOR2_X1 U25077 ( .A1(n11382), .A2(n2756), .ZN(n2819) );
NOR2_X1 U25078 ( .A1(n11379), .A2(n2756), .ZN(n2778) );
NOR2_X1 U25079 ( .A1(n11377), .A2(n2756), .ZN(n2785) );
NOR2_X1 U25080 ( .A1(n11375), .A2(n2756), .ZN(n2866) );
NOR2_X1 U25081 ( .A1(n11380), .A2(n2756), .ZN(n2808) );
NOR2_X1 U25082 ( .A1(n11378), .A2(n2756), .ZN(n2791) );
NOR2_X1 U25083 ( .A1(n11384), .A2(n2756), .ZN(n2825) );
NOR2_X1 U25084 ( .A1(n11385), .A2(n2756), .ZN(n2854) );
NAND2_X1 U25085 ( .A1(n2871), .A2(n2872), .ZN(n2437) );
NOR2_X1 U25086 ( .A1(n2876), .A2(n2877), .ZN(n2871) );
NOR2_X1 U25087 ( .A1(n2873), .A2(n2874), .ZN(n2872) );
NOR2_X1 U25088 ( .A1(n11371), .A2(n2169), .ZN(n2876) );
NAND2_X1 U25089 ( .A1(n2783), .A2(n2784), .ZN(n2043) );
NOR2_X1 U25090 ( .A1(n2787), .A2(n2788), .ZN(n2783) );
NOR2_X1 U25091 ( .A1(n2785), .A2(n2786), .ZN(n2784) );
NOR2_X1 U25092 ( .A1(n11349), .A2(n16448), .ZN(n2787) );
NAND2_X1 U25093 ( .A1(n11318), .A2(n11504), .ZN(n10377) );
NOR2_X1 U25094 ( .A1(n10148), .A2(n10149), .ZN(n10146) );
NOR2_X1 U25095 ( .A1(n10150), .A2(n11328), .ZN(n10149) );
NAND2_X1 U25096 ( .A1(n10459), .A2(n10545), .ZN(n5182) );
AND2_X1 U25097 ( .A1(n10547), .A2(n10546), .ZN(n10459) );
NAND2_X1 U25098 ( .A1(n11312), .A2(n15810), .ZN(n10173) );
NAND2_X1 U25099 ( .A1(n10470), .A2(n10471), .ZN(n5162) );
NOR2_X1 U25100 ( .A1(n15819), .A2(n15800), .ZN(n10470) );
NOR2_X1 U25101 ( .A1(n11516), .A2(n15798), .ZN(n10471) );
NAND2_X1 U25102 ( .A1(n11498), .A2(n5217), .ZN(n5151) );
NAND2_X1 U25103 ( .A1(n5218), .A2(n5131), .ZN(n5217) );
NOR2_X1 U25104 ( .A1(debug_req_i), .A2(n5133), .ZN(n5218) );
NAND2_X1 U25105 ( .A1(n3594), .A2(n3595), .ZN(n1449) );
NAND2_X1 U25106 ( .A1(n3596), .A2(n2863), .ZN(n3595) );
NAND2_X1 U25107 ( .A1(n3599), .A2(n3600), .ZN(n3596) );
NAND2_X1 U25108 ( .A1(instr_rdata_i_16_), .A2(n11460), .ZN(n3600) );
NAND2_X1 U25109 ( .A1(n2823), .A2(n2824), .ZN(n2308) );
NOR2_X1 U25110 ( .A1(n2827), .A2(n2828), .ZN(n2823) );
NOR2_X1 U25111 ( .A1(n2825), .A2(n2826), .ZN(n2824) );
NOR2_X1 U25112 ( .A1(n11363), .A2(n2169), .ZN(n2827) );
NAND2_X1 U25113 ( .A1(n10543), .A2(n10544), .ZN(n10144) );
NOR2_X1 U25114 ( .A1(n15799), .A2(n15814), .ZN(n10543) );
NOR2_X1 U25115 ( .A1(n11326), .A2(n10523), .ZN(n10544) );
INV_X1 U25116 ( .A(instr_rdata_i_0_), .ZN(n19961) );
INV_X1 U25117 ( .A(instr_rdata_i_16_), .ZN(n19945) );
NOR2_X1 U25118 ( .A1(n10525), .A2(n10233), .ZN(n10524) );
OR2_X1 U25119 ( .A1(n11327), .A2(n10523), .ZN(n10525) );
NAND2_X1 U25120 ( .A1(n10309), .A2(n10310), .ZN(n5167) );
NOR2_X1 U25121 ( .A1(n15798), .A2(n15915), .ZN(n10309) );
NOR2_X1 U25122 ( .A1(n11514), .A2(n11517), .ZN(n10310) );
INV_X1 U25123 ( .A(instr_rdata_i_12_), .ZN(n19949) );
INV_X1 U25124 ( .A(instr_rdata_i_11_), .ZN(n19950) );
INV_X1 U25125 ( .A(instr_rdata_i_10_), .ZN(n19951) );
INV_X1 U25126 ( .A(instr_rdata_i_7_), .ZN(n19954) );
INV_X1 U25127 ( .A(instr_rdata_i_4_), .ZN(n19957) );
INV_X1 U25128 ( .A(instr_rdata_i_2_), .ZN(n19959) );
INV_X1 U25129 ( .A(instr_rdata_i_31_), .ZN(n19908) );
INV_X1 U25130 ( .A(instr_rdata_i_28_), .ZN(n19915) );
INV_X1 U25131 ( .A(instr_rdata_i_27_), .ZN(n19918) );
INV_X1 U25132 ( .A(instr_rdata_i_26_), .ZN(n19920) );
INV_X1 U25133 ( .A(instr_rdata_i_23_), .ZN(n19926) );
INV_X1 U25134 ( .A(instr_rdata_i_20_), .ZN(n19932) );
INV_X1 U25135 ( .A(instr_rdata_i_18_), .ZN(n19935) );
INV_X1 U25136 ( .A(instr_rdata_i_15_), .ZN(n19946) );
INV_X1 U25137 ( .A(instr_rdata_i_9_), .ZN(n19952) );
NAND2_X1 U25138 ( .A1(n10461), .A2(n11517), .ZN(n5142) );
NOR2_X1 U25139 ( .A1(n11401), .A2(n2164), .ZN(n2633) );
NOR2_X1 U25140 ( .A1(n11403), .A2(n2164), .ZN(n2576) );
NOR2_X1 U25141 ( .A1(n11402), .A2(n2164), .ZN(n2605) );
NOR2_X1 U25142 ( .A1(n11398), .A2(n2164), .ZN(n2163) );
NOR2_X1 U25143 ( .A1(n11393), .A2(n2164), .ZN(n2284) );
NOR2_X1 U25144 ( .A1(n11424), .A2(n2164), .ZN(n2327) );
NOR2_X1 U25145 ( .A1(n10608), .A2(n16444), .ZN(n2937) );
NOR2_X1 U25146 ( .A1(n10606), .A2(n16444), .ZN(n2925) );
NOR2_X1 U25147 ( .A1(n10604), .A2(n2900), .ZN(n2921) );
NOR2_X1 U25148 ( .A1(n10602), .A2(n2900), .ZN(n2917) );
NOR2_X1 U25149 ( .A1(n10600), .A2(n2900), .ZN(n2913) );
NOR2_X1 U25150 ( .A1(n10598), .A2(n16444), .ZN(n2909) );
NOR2_X1 U25151 ( .A1(n10596), .A2(n2900), .ZN(n2905) );
NOR2_X1 U25152 ( .A1(n10594), .A2(n16444), .ZN(n2899) );
NOR2_X1 U25153 ( .A1(n10592), .A2(n16444), .ZN(n3017) );
NOR2_X1 U25154 ( .A1(n10588), .A2(n2900), .ZN(n3009) );
NOR2_X1 U25155 ( .A1(n10586), .A2(n16444), .ZN(n3005) );
NOR2_X1 U25156 ( .A1(n10584), .A2(n2900), .ZN(n3001) );
NOR2_X1 U25157 ( .A1(n10582), .A2(n2900), .ZN(n2997) );
NOR2_X1 U25158 ( .A1(n10578), .A2(n16444), .ZN(n2989) );
NOR2_X1 U25159 ( .A1(n10576), .A2(n2900), .ZN(n2985) );
NOR2_X1 U25160 ( .A1(n10574), .A2(n2900), .ZN(n2981) );
NOR2_X1 U25161 ( .A1(n10570), .A2(n16444), .ZN(n2973) );
NOR2_X1 U25162 ( .A1(n10568), .A2(n16444), .ZN(n2969) );
NOR2_X1 U25163 ( .A1(n10566), .A2(n2900), .ZN(n2965) );
NOR2_X1 U25164 ( .A1(n10564), .A2(n16444), .ZN(n2961) );
NOR2_X1 U25165 ( .A1(n10560), .A2(n2900), .ZN(n2953) );
NOR2_X1 U25166 ( .A1(n10554), .A2(n2900), .ZN(n2941) );
NOR2_X1 U25167 ( .A1(n10552), .A2(n2900), .ZN(n2933) );
NOR2_X1 U25168 ( .A1(n10550), .A2(n16444), .ZN(n2929) );
NOR2_X1 U25169 ( .A1(n10644), .A2(n20927), .ZN(n3501) );
NOR2_X1 U25170 ( .A1(n2187), .A2(n2117), .ZN(n2185) );
NOR2_X1 U25171 ( .A1(n2188), .A2(n2189), .ZN(n2187) );
NAND2_X1 U25172 ( .A1(n2190), .A2(n2191), .ZN(n2189) );
NOR2_X1 U25173 ( .A1(n11381), .A2(n2169), .ZN(n2188) );
NOR2_X1 U25174 ( .A1(n10725), .A2(n20927), .ZN(n4007) );
NOR2_X1 U25175 ( .A1(n10753), .A2(n20927), .ZN(n3982) );
NOR2_X1 U25176 ( .A1(n10768), .A2(n20927), .ZN(n3959) );
NOR2_X1 U25177 ( .A1(n10787), .A2(n20927), .ZN(n3948) );
NOR2_X1 U25178 ( .A1(n10802), .A2(n20927), .ZN(n3937) );
NOR2_X1 U25179 ( .A1(n10816), .A2(n20927), .ZN(n3926) );
NOR2_X1 U25180 ( .A1(n10646), .A2(n20927), .ZN(n3903) );
NOR2_X1 U25181 ( .A1(n10846), .A2(n20927), .ZN(n3892) );
NOR2_X1 U25182 ( .A1(n10863), .A2(n20927), .ZN(n3881) );
NOR2_X1 U25183 ( .A1(n10617), .A2(n20927), .ZN(n3858) );
NOR2_X1 U25184 ( .A1(n10893), .A2(n20927), .ZN(n3847) );
NOR2_X1 U25185 ( .A1(n10908), .A2(n20927), .ZN(n3836) );
NOR2_X1 U25186 ( .A1(n10923), .A2(n20927), .ZN(n3825) );
NOR2_X1 U25187 ( .A1(n10953), .A2(n20927), .ZN(n3802) );
NOR2_X1 U25188 ( .A1(n10661), .A2(n20927), .ZN(n3728) );
NOR2_X1 U25189 ( .A1(n10669), .A2(n20927), .ZN(n4057) );
NOR2_X1 U25190 ( .A1(n10698), .A2(n20927), .ZN(n4038) );
NOR2_X1 U25191 ( .A1(n10711), .A2(n20927), .ZN(n4022) );
NOR2_X1 U25192 ( .A1(n10621), .A2(n20927), .ZN(n3763) );
NOR2_X1 U25193 ( .A1(n10615), .A2(n20927), .ZN(n3752) );
NOR2_X1 U25194 ( .A1(n10610), .A2(n20927), .ZN(n4030) );
NOR2_X1 U25195 ( .A1(n10679), .A2(n20927), .ZN(n4014) );
NOR2_X1 U25196 ( .A1(n10739), .A2(n20927), .ZN(n3993) );
NOR2_X1 U25197 ( .A1(n10981), .A2(n20927), .ZN(n3741) );
NOR2_X1 U25198 ( .A1(n11007), .A2(n16354), .ZN(n7572) );
NOR2_X1 U25199 ( .A1(n10980), .A2(n20924), .ZN(n7374) );
NOR2_X1 U25200 ( .A1(n10978), .A2(n20924), .ZN(n7550) );
NOR2_X1 U25201 ( .A1(n10967), .A2(n20924), .ZN(n7414) );
NOR2_X1 U25202 ( .A1(n10952), .A2(n20924), .ZN(n7422) );
NOR2_X1 U25203 ( .A1(n10937), .A2(n20924), .ZN(n7430) );
NOR2_X1 U25204 ( .A1(n10922), .A2(n20924), .ZN(n7438) );
NOR2_X1 U25205 ( .A1(n10907), .A2(n20924), .ZN(n7446) );
NOR2_X1 U25206 ( .A1(n10892), .A2(n20924), .ZN(n7454) );
NOR2_X1 U25207 ( .A1(n10877), .A2(n16354), .ZN(n7470) );
NOR2_X1 U25208 ( .A1(n10862), .A2(n16354), .ZN(n7486) );
NOR2_X1 U25209 ( .A1(n10845), .A2(n20924), .ZN(n7494) );
NOR2_X1 U25210 ( .A1(n10830), .A2(n16354), .ZN(n7510) );
NOR2_X1 U25211 ( .A1(n10815), .A2(n16354), .ZN(n7518) );
NOR2_X1 U25212 ( .A1(n10801), .A2(n16354), .ZN(n7526) );
NOR2_X1 U25213 ( .A1(n10786), .A2(n20924), .ZN(n7534) );
NOR2_X1 U25214 ( .A1(n10767), .A2(n20924), .ZN(n7542) );
NOR2_X1 U25215 ( .A1(n10752), .A2(n20924), .ZN(n7558) );
NOR2_X1 U25216 ( .A1(n10724), .A2(n20924), .ZN(n7326) );
NOR2_X1 U25217 ( .A1(n10710), .A2(n16354), .ZN(n7342) );
NOR2_X1 U25218 ( .A1(n10697), .A2(n16354), .ZN(n7358) );
NOR2_X1 U25219 ( .A1(n10678), .A2(n20924), .ZN(n7334) );
NOR2_X1 U25220 ( .A1(n10668), .A2(n16354), .ZN(n7366) );
NOR2_X1 U25221 ( .A1(n10660), .A2(n16354), .ZN(n7390) );
NOR2_X1 U25222 ( .A1(n10645), .A2(n20924), .ZN(n7502) );
NOR2_X1 U25223 ( .A1(n10643), .A2(n16354), .ZN(n7478) );
NOR2_X1 U25224 ( .A1(n10630), .A2(n16354), .ZN(n7406) );
NOR2_X1 U25225 ( .A1(n10620), .A2(n16354), .ZN(n7398) );
NOR2_X1 U25226 ( .A1(n10616), .A2(n16354), .ZN(n7462) );
NOR2_X1 U25227 ( .A1(n10614), .A2(n20924), .ZN(n7382) );
NOR2_X1 U25228 ( .A1(n10609), .A2(n20924), .ZN(n7350) );
NOR2_X1 U25229 ( .A1(n11384), .A2(n16448), .ZN(n2659) );
NOR2_X1 U25230 ( .A1(n11462), .A2(n16448), .ZN(n2636) );
NOR2_X1 U25231 ( .A1(n11031), .A2(n16365), .ZN(n9427) );
NOR2_X1 U25232 ( .A1(n11033), .A2(n16365), .ZN(n8870) );
NOR2_X1 U25233 ( .A1(n11034), .A2(n16365), .ZN(n8818) );
NOR2_X1 U25234 ( .A1(n11382), .A2(n16448), .ZN(n2168) );
NOR2_X1 U25235 ( .A1(n11377), .A2(n2169), .ZN(n2287) );
NOR2_X1 U25236 ( .A1(n11375), .A2(n2169), .ZN(n2330) );
NOR2_X1 U25237 ( .A1(n2249), .A2(n2117), .ZN(n2248) );
NOR2_X1 U25238 ( .A1(n2250), .A2(n2251), .ZN(n2249) );
NAND2_X1 U25239 ( .A1(n2252), .A2(n2253), .ZN(n2251) );
NOR2_X1 U25240 ( .A1(n11378), .A2(n2169), .ZN(n2250) );
INV_X1 U25241 ( .A(data_gnt_i), .ZN(n19965) );
NOR2_X1 U25242 ( .A1(n10662), .A2(n8773), .ZN(n9888) );
NOR2_X1 U25243 ( .A1(n11465), .A2(n8773), .ZN(n9425) );
NOR2_X1 U25244 ( .A1(n10670), .A2(n8773), .ZN(n8868) );
NOR2_X1 U25245 ( .A1(n10704), .A2(n8773), .ZN(n8816) );
NAND2_X1 U25246 ( .A1(n6543), .A2(n20938), .ZN(n6540) );
AND2_X1 U25247 ( .A1(n6545), .A2(n11320), .ZN(n6543) );
NAND2_X1 U25248 ( .A1(n11332), .A2(n10390), .ZN(n5258) );
NAND2_X1 U25249 ( .A1(n21534), .A2(crash_dump_o_110_), .ZN(n21540) );
NOR2_X1 U25250 ( .A1(n21533), .A2(n10788), .ZN(n21534) );
NAND2_X1 U25251 ( .A1(n21541), .A2(crash_dump_o_112_), .ZN(n21547) );
NOR2_X1 U25252 ( .A1(n21540), .A2(n10817), .ZN(n21541) );
NAND2_X1 U25253 ( .A1(n21548), .A2(crash_dump_o_114_), .ZN(n21556) );
NOR2_X1 U25254 ( .A1(n21547), .A2(n10647), .ZN(n21548) );
NAND2_X1 U25255 ( .A1(n21557), .A2(crash_dump_o_116_), .ZN(n21563) );
NOR2_X1 U25256 ( .A1(n21556), .A2(n10864), .ZN(n21557) );
NAND2_X1 U25257 ( .A1(n21564), .A2(crash_dump_o_118_), .ZN(n21570) );
NOR2_X1 U25258 ( .A1(n21563), .A2(n11495), .ZN(n21564) );
NAND2_X1 U25259 ( .A1(n21571), .A2(crash_dump_o_120_), .ZN(n21577) );
NOR2_X1 U25260 ( .A1(n21570), .A2(n10909), .ZN(n21571) );
NAND2_X1 U25261 ( .A1(n21578), .A2(crash_dump_o_122_), .ZN(n21584) );
NOR2_X1 U25262 ( .A1(n21577), .A2(n10939), .ZN(n21578) );
NAND2_X1 U25263 ( .A1(n22514), .A2(cs_registers_i_mhpmcounter_2__58_), .ZN(n22522) );
NOR2_X1 U25264 ( .A1(n22513), .A2(n10936), .ZN(n22514) );
NAND2_X1 U25265 ( .A1(n22417), .A2(cs_registers_i_mhpmcounter_2__32_), .ZN(n22423) );
NOR2_X1 U25266 ( .A1(n22416), .A2(n11126), .ZN(n22417) );
NAND2_X1 U25267 ( .A1(n22410), .A2(cs_registers_i_mhpmcounter_2__30_), .ZN(n22416) );
NOR2_X1 U25268 ( .A1(n22409), .A2(n11491), .ZN(n22410) );
NAND2_X1 U25269 ( .A1(n22400), .A2(cs_registers_i_mhpmcounter_2__28_), .ZN(n22409) );
NOR2_X1 U25270 ( .A1(n22399), .A2(n10965), .ZN(n22400) );
NAND2_X1 U25271 ( .A1(n22199), .A2(cs_registers_i_mhpmcounter_0__32_), .ZN(n22205) );
NOR2_X1 U25272 ( .A1(n22198), .A2(n11510), .ZN(n22199) );
NAND2_X1 U25273 ( .A1(n22192), .A2(cs_registers_i_mhpmcounter_0__30_), .ZN(n22198) );
NOR2_X1 U25274 ( .A1(n22191), .A2(n10625), .ZN(n22192) );
NAND2_X1 U25275 ( .A1(n22182), .A2(cs_registers_i_mhpmcounter_0__28_), .ZN(n22191) );
NOR2_X1 U25276 ( .A1(n22181), .A2(n10963), .ZN(n22182) );
NAND2_X1 U25277 ( .A1(n21520), .A2(crash_dump_o_106_), .ZN(n21526) );
NOR2_X1 U25278 ( .A1(n10745), .A2(n21616), .ZN(n21520) );
NAND2_X1 U25279 ( .A1(n21465), .A2(crash_dump_o_88_), .ZN(n21471) );
NOR2_X1 U25280 ( .A1(n21464), .A2(n10910), .ZN(n21465) );
NAND2_X1 U25281 ( .A1(n22507), .A2(cs_registers_i_mhpmcounter_2__56_), .ZN(n22513) );
NOR2_X1 U25282 ( .A1(n22506), .A2(n10906), .ZN(n22507) );
NAND2_X1 U25283 ( .A1(n22386), .A2(cs_registers_i_mhpmcounter_2__24_), .ZN(n22392) );
NOR2_X1 U25284 ( .A1(n22385), .A2(n10905), .ZN(n22386) );
NAND2_X1 U25285 ( .A1(n22289), .A2(cs_registers_i_mhpmcounter_0__56_), .ZN(n22295) );
NOR2_X1 U25286 ( .A1(n22288), .A2(n10904), .ZN(n22289) );
NAND2_X1 U25287 ( .A1(n22168), .A2(cs_registers_i_mhpmcounter_0__24_), .ZN(n22174) );
NOR2_X1 U25288 ( .A1(n22167), .A2(n10903), .ZN(n22168) );
NAND2_X1 U25289 ( .A1(n21458), .A2(crash_dump_o_86_), .ZN(n21464) );
NOR2_X1 U25290 ( .A1(n21457), .A2(n11496), .ZN(n21458) );
NAND2_X1 U25291 ( .A1(n22500), .A2(cs_registers_i_mhpmcounter_2__54_), .ZN(n22506) );
NOR2_X1 U25292 ( .A1(n22499), .A2(n11131), .ZN(n22500) );
NAND2_X1 U25293 ( .A1(n22379), .A2(cs_registers_i_mhpmcounter_2__22_), .ZN(n22385) );
NOR2_X1 U25294 ( .A1(n22378), .A2(n11123), .ZN(n22379) );
NAND2_X1 U25295 ( .A1(n22282), .A2(cs_registers_i_mhpmcounter_0__54_), .ZN(n22288) );
NOR2_X1 U25296 ( .A1(n22281), .A2(n11120), .ZN(n22282) );
NAND2_X1 U25297 ( .A1(n22161), .A2(cs_registers_i_mhpmcounter_0__22_), .ZN(n22167) );
NOR2_X1 U25298 ( .A1(n22160), .A2(n11114), .ZN(n22161) );
NAND2_X1 U25299 ( .A1(n21451), .A2(crash_dump_o_84_), .ZN(n21457) );
NOR2_X1 U25300 ( .A1(n21450), .A2(n10865), .ZN(n21451) );
NAND2_X1 U25301 ( .A1(n22493), .A2(cs_registers_i_mhpmcounter_2__52_), .ZN(n22499) );
NOR2_X1 U25302 ( .A1(n22492), .A2(n10861), .ZN(n22493) );
NAND2_X1 U25303 ( .A1(n22372), .A2(cs_registers_i_mhpmcounter_2__20_), .ZN(n22378) );
NOR2_X1 U25304 ( .A1(n22371), .A2(n10860), .ZN(n22372) );
NAND2_X1 U25305 ( .A1(n22275), .A2(cs_registers_i_mhpmcounter_0__52_), .ZN(n22281) );
NOR2_X1 U25306 ( .A1(n22274), .A2(n10859), .ZN(n22275) );
NAND2_X1 U25307 ( .A1(n22154), .A2(cs_registers_i_mhpmcounter_0__20_), .ZN(n22160) );
NOR2_X1 U25308 ( .A1(n22153), .A2(n10858), .ZN(n22154) );
NAND2_X1 U25309 ( .A1(n21438), .A2(crash_dump_o_82_), .ZN(n21450) );
NOR2_X1 U25310 ( .A1(n21437), .A2(n10648), .ZN(n21438) );
NAND2_X1 U25311 ( .A1(n22486), .A2(cs_registers_i_mhpmcounter_2__50_), .ZN(n22492) );
NOR2_X1 U25312 ( .A1(n22485), .A2(n10653), .ZN(n22486) );
NAND2_X1 U25313 ( .A1(n22363), .A2(cs_registers_i_mhpmcounter_2__18_), .ZN(n22371) );
NOR2_X1 U25314 ( .A1(n22362), .A2(n10652), .ZN(n22363) );
NAND2_X1 U25315 ( .A1(n22268), .A2(cs_registers_i_mhpmcounter_0__50_), .ZN(n22274) );
NOR2_X1 U25316 ( .A1(n22267), .A2(n10651), .ZN(n22268) );
NAND2_X1 U25317 ( .A1(n22145), .A2(cs_registers_i_mhpmcounter_0__18_), .ZN(n22153) );
NOR2_X1 U25318 ( .A1(n22144), .A2(n10650), .ZN(n22145) );
NAND2_X1 U25319 ( .A1(n21431), .A2(crash_dump_o_80_), .ZN(n21437) );
NOR2_X1 U25320 ( .A1(n21430), .A2(n10818), .ZN(n21431) );
NAND2_X1 U25321 ( .A1(n22475), .A2(cs_registers_i_mhpmcounter_2__48_), .ZN(n22485) );
NOR2_X1 U25322 ( .A1(n22474), .A2(n10814), .ZN(n22475) );
NAND2_X1 U25323 ( .A1(n22356), .A2(cs_registers_i_mhpmcounter_2__16_), .ZN(n22362) );
NOR2_X1 U25324 ( .A1(n22355), .A2(n10813), .ZN(n22356) );
NAND2_X1 U25325 ( .A1(n22257), .A2(cs_registers_i_mhpmcounter_0__48_), .ZN(n22267) );
NOR2_X1 U25326 ( .A1(n22256), .A2(n10812), .ZN(n22257) );
NAND2_X1 U25327 ( .A1(n22138), .A2(cs_registers_i_mhpmcounter_0__16_), .ZN(n22144) );
NOR2_X1 U25328 ( .A1(n22137), .A2(n10811), .ZN(n22138) );
NAND2_X1 U25329 ( .A1(n21424), .A2(crash_dump_o_78_), .ZN(n21430) );
NOR2_X1 U25330 ( .A1(n21423), .A2(n10789), .ZN(n21424) );
NAND2_X1 U25331 ( .A1(n22468), .A2(cs_registers_i_mhpmcounter_2__46_), .ZN(n22474) );
NOR2_X1 U25332 ( .A1(n22467), .A2(n10785), .ZN(n22468) );
NAND2_X1 U25333 ( .A1(n22349), .A2(cs_registers_i_mhpmcounter_2__14_), .ZN(n22355) );
NOR2_X1 U25334 ( .A1(n22348), .A2(n10784), .ZN(n22349) );
NAND2_X1 U25335 ( .A1(n22250), .A2(cs_registers_i_mhpmcounter_0__46_), .ZN(n22256) );
NOR2_X1 U25336 ( .A1(n22249), .A2(n10783), .ZN(n22250) );
NAND2_X1 U25337 ( .A1(n22131), .A2(cs_registers_i_mhpmcounter_0__14_), .ZN(n22137) );
NOR2_X1 U25338 ( .A1(n22130), .A2(n10782), .ZN(n22131) );
NAND2_X1 U25339 ( .A1(n21527), .A2(crash_dump_o_108_), .ZN(n21533) );
NOR2_X1 U25340 ( .A1(n21526), .A2(n11307), .ZN(n21527) );
NAND2_X1 U25341 ( .A1(n21417), .A2(crash_dump_o_76_), .ZN(n21423) );
NOR2_X1 U25342 ( .A1(n21416), .A2(n11308), .ZN(n21417) );
NAND2_X1 U25343 ( .A1(n22461), .A2(cs_registers_i_mhpmcounter_2__44_), .ZN(n22467) );
NOR2_X1 U25344 ( .A1(n22460), .A2(n10764), .ZN(n22461) );
NAND2_X1 U25345 ( .A1(n22342), .A2(cs_registers_i_mhpmcounter_2__12_), .ZN(n22348) );
NOR2_X1 U25346 ( .A1(n22341), .A2(n10763), .ZN(n22342) );
NAND2_X1 U25347 ( .A1(n22243), .A2(cs_registers_i_mhpmcounter_0__44_), .ZN(n22249) );
NOR2_X1 U25348 ( .A1(n22242), .A2(n10762), .ZN(n22243) );
NAND2_X1 U25349 ( .A1(n22124), .A2(cs_registers_i_mhpmcounter_0__12_), .ZN(n22130) );
NOR2_X1 U25350 ( .A1(n22123), .A2(n10761), .ZN(n22124) );
NAND2_X1 U25351 ( .A1(n22454), .A2(cs_registers_i_mhpmcounter_2__42_), .ZN(n22460) );
NOR2_X1 U25352 ( .A1(n22453), .A2(n10735), .ZN(n22454) );
NAND2_X1 U25353 ( .A1(n22335), .A2(cs_registers_i_mhpmcounter_2__10_), .ZN(n22341) );
NOR2_X1 U25354 ( .A1(n10736), .A2(n22543), .ZN(n22335) );
NAND2_X1 U25355 ( .A1(n22236), .A2(cs_registers_i_mhpmcounter_0__42_), .ZN(n22242) );
NOR2_X1 U25356 ( .A1(n22235), .A2(n10733), .ZN(n22236) );
NAND2_X1 U25357 ( .A1(n22117), .A2(cs_registers_i_mhpmcounter_0__10_), .ZN(n22123) );
NOR2_X1 U25358 ( .A1(n10734), .A2(n22325), .ZN(n22117) );
NAND2_X1 U25359 ( .A1(n21410), .A2(crash_dump_o_74_), .ZN(n21416) );
NOR2_X1 U25360 ( .A1(n21509), .A2(n10746), .ZN(n21410) );
NAND2_X1 U25361 ( .A1(n21409), .A2(crash_dump_o_72_), .ZN(n21509) );
NOR2_X1 U25362 ( .A1(n21503), .A2(n10681), .ZN(n21409) );
NAND2_X1 U25363 ( .A1(n22447), .A2(cs_registers_i_mhpmcounter_2__40_), .ZN(n22453) );
NOR2_X1 U25364 ( .A1(n22446), .A2(n10685), .ZN(n22447) );
NAND2_X1 U25365 ( .A1(n22229), .A2(cs_registers_i_mhpmcounter_0__40_), .ZN(n22235) );
NOR2_X1 U25366 ( .A1(n22228), .A2(n10683), .ZN(n22229) );
NAND2_X1 U25367 ( .A1(n21408), .A2(crash_dump_o_70_), .ZN(n21503) );
NOR2_X1 U25368 ( .A1(n21497), .A2(n11513), .ZN(n21408) );
NAND2_X1 U25369 ( .A1(n21515), .A2(crash_dump_o_102_), .ZN(n21612) );
NOR2_X1 U25370 ( .A1(n21606), .A2(n11466), .ZN(n21515) );
NAND2_X1 U25371 ( .A1(n22330), .A2(cs_registers_i_mhpmcounter_2__6_), .ZN(n22539) );
NOR2_X1 U25372 ( .A1(n22533), .A2(n11132), .ZN(n22330) );
NAND2_X1 U25373 ( .A1(n22438), .A2(cs_registers_i_mhpmcounter_2__38_), .ZN(n22446) );
NOR2_X1 U25374 ( .A1(n22437), .A2(n11130), .ZN(n22438) );
NAND2_X1 U25375 ( .A1(n22112), .A2(cs_registers_i_mhpmcounter_0__6_), .ZN(n22321) );
NOR2_X1 U25376 ( .A1(n22315), .A2(n11121), .ZN(n22112) );
NAND2_X1 U25377 ( .A1(n22220), .A2(cs_registers_i_mhpmcounter_0__38_), .ZN(n22228) );
NOR2_X1 U25378 ( .A1(n22219), .A2(n11119), .ZN(n22220) );
NAND2_X1 U25379 ( .A1(n22431), .A2(cs_registers_i_mhpmcounter_2__36_), .ZN(n22437) );
NOR2_X1 U25380 ( .A1(n22430), .A2(n10674), .ZN(n22431) );
NAND2_X1 U25381 ( .A1(n22213), .A2(cs_registers_i_mhpmcounter_0__36_), .ZN(n22219) );
NOR2_X1 U25382 ( .A1(n22212), .A2(n10673), .ZN(n22213) );
NAND2_X1 U25383 ( .A1(n22328), .A2(cs_registers_i_mhpmcounter_2__2_), .ZN(n22478) );
NOR2_X1 U25384 ( .A1(n11479), .A2(n11122), .ZN(n22328) );
NAND2_X1 U25385 ( .A1(n22424), .A2(cs_registers_i_mhpmcounter_2__34_), .ZN(n22430) );
NOR2_X1 U25386 ( .A1(n22423), .A2(n11128), .ZN(n22424) );
NAND2_X1 U25387 ( .A1(n22206), .A2(cs_registers_i_mhpmcounter_0__34_), .ZN(n22212) );
NOR2_X1 U25388 ( .A1(n22205), .A2(n11117), .ZN(n22206) );
NAND2_X1 U25389 ( .A1(n22393), .A2(cs_registers_i_mhpmcounter_2__26_), .ZN(n22399) );
NOR2_X1 U25390 ( .A1(n22392), .A2(n10935), .ZN(n22393) );
NAND2_X1 U25391 ( .A1(n22296), .A2(cs_registers_i_mhpmcounter_0__58_), .ZN(n22304) );
NOR2_X1 U25392 ( .A1(n22295), .A2(n10934), .ZN(n22296) );
NAND2_X1 U25393 ( .A1(n22175), .A2(cs_registers_i_mhpmcounter_0__26_), .ZN(n22181) );
NOR2_X1 U25394 ( .A1(n22174), .A2(n10933), .ZN(n22175) );
NAND2_X1 U25395 ( .A1(n21472), .A2(crash_dump_o_90_), .ZN(n21478) );
NOR2_X1 U25396 ( .A1(n21471), .A2(n10940), .ZN(n21472) );
NAND2_X1 U25397 ( .A1(n21486), .A2(crash_dump_o_68_), .ZN(n21497) );
NAND2_X1 U25398 ( .A1(n22110), .A2(cs_registers_i_mhpmcounter_0__2_), .ZN(n22260) );
NOR2_X1 U25399 ( .A1(n10665), .A2(n10666), .ZN(n22110) );
NAND2_X1 U25400 ( .A1(n22329), .A2(cs_registers_i_mhpmcounter_2__4_), .ZN(n22533) );
NOR2_X1 U25401 ( .A1(n22478), .A2(n10675), .ZN(n22329) );
NAND2_X1 U25402 ( .A1(n22111), .A2(cs_registers_i_mhpmcounter_0__4_), .ZN(n22315) );
NOR2_X1 U25403 ( .A1(n22260), .A2(n11478), .ZN(n22111) );
NAND2_X1 U25404 ( .A1(n21514), .A2(crash_dump_o_100_), .ZN(n21606) );
NOR2_X1 U25405 ( .A1(n21600), .A2(n10670), .ZN(n21514) );
NAND2_X1 U25406 ( .A1(n21513), .A2(instr_fetch_err_plus2), .ZN(n21600) );
NOR2_X1 U25407 ( .A1(n11465), .A2(n10662), .ZN(n21513) );
NAND2_X1 U25408 ( .A1(n11326), .A2(n15799), .ZN(n10233) );
NOR2_X1 U25409 ( .A1(n11467), .A2(n16392), .ZN(n7378) );
NOR2_X1 U25410 ( .A1(n10745), .A2(n16392), .ZN(n7320) );
NOR2_X1 U25411 ( .A1(n10731), .A2(n16392), .ZN(n7330) );
NOR2_X1 U25412 ( .A1(n10717), .A2(n16392), .ZN(n7346) );
NOR2_X1 U25413 ( .A1(n10704), .A2(n16392), .ZN(n7362) );
NOR2_X1 U25414 ( .A1(n10680), .A2(n16392), .ZN(n7338) );
NOR2_X1 U25415 ( .A1(n10670), .A2(n16392), .ZN(n7370) );
NOR2_X1 U25416 ( .A1(n11466), .A2(n16392), .ZN(n7354) );
NOR2_X1 U25417 ( .A1(n11185), .A2(n16419), .ZN(n4898) );
NOR2_X1 U25418 ( .A1(n11187), .A2(n16419), .ZN(n4879) );
NOR2_X1 U25419 ( .A1(n11188), .A2(n16419), .ZN(n4860) );
NOR2_X1 U25420 ( .A1(n11189), .A2(n16419), .ZN(n4841) );
NOR2_X1 U25421 ( .A1(n11190), .A2(n16419), .ZN(n4822) );
NOR2_X1 U25422 ( .A1(n11191), .A2(n16419), .ZN(n4803) );
NOR2_X1 U25423 ( .A1(n11192), .A2(n16419), .ZN(n4781) );
NOR2_X1 U25424 ( .A1(n11193), .A2(n16419), .ZN(n4760) );
NAND2_X1 U25425 ( .A1(n21516), .A2(crash_dump_o_104_), .ZN(n21616) );
NOR2_X1 U25426 ( .A1(n21612), .A2(n10680), .ZN(n21516) );
NAND2_X1 U25427 ( .A1(n22331), .A2(cs_registers_i_mhpmcounter_2__8_), .ZN(n22543) );
NOR2_X1 U25428 ( .A1(n22539), .A2(n10686), .ZN(n22331) );
NAND2_X1 U25429 ( .A1(n22113), .A2(cs_registers_i_mhpmcounter_0__8_), .ZN(n22325) );
NOR2_X1 U25430 ( .A1(n22321), .A2(n10684), .ZN(n22113) );
NAND2_X1 U25431 ( .A1(n10452), .A2(n10453), .ZN(n10070) );
NOR2_X1 U25432 ( .A1(n11502), .A2(n11504), .ZN(n10453) );
NOR2_X1 U25433 ( .A1(n15884), .A2(n1440), .ZN(n10452) );
NAND2_X1 U25434 ( .A1(n11333), .A2(n11328), .ZN(n5580) );
NAND2_X1 U25435 ( .A1(n11338), .A2(n10390), .ZN(n10286) );
NAND2_X1 U25436 ( .A1(n11298), .A2(n1579), .ZN(n1575) );
NAND2_X1 U25437 ( .A1(n10264), .A2(n10265), .ZN(n10097) );
NOR2_X1 U25438 ( .A1(n15914), .A2(n15816), .ZN(n10264) );
NOR2_X1 U25439 ( .A1(n11328), .A2(n15860), .ZN(n10265) );
NAND2_X1 U25440 ( .A1(n11062), .A2(n15822), .ZN(n1304) );
NAND2_X1 U25441 ( .A1(n11322), .A2(n11326), .ZN(n10244) );
NAND2_X1 U25442 ( .A1(n10539), .A2(n11298), .ZN(n1554) );
NOR2_X1 U25443 ( .A1(n11295), .A2(n15825), .ZN(n10539) );
NAND2_X1 U25444 ( .A1(instr_gnt_i), .A2(instr_req_o), .ZN(n3028) );
NAND2_X1 U25445 ( .A1(n10439), .A2(n11311), .ZN(n10433) );
NOR2_X1 U25446 ( .A1(n15807), .A2(n15892), .ZN(n10439) );
NAND2_X1 U25447 ( .A1(n11312), .A2(n11319), .ZN(n10188) );
NOR2_X1 U25448 ( .A1(n11513), .A2(n16389), .ZN(n7897) );
NOR2_X1 U25449 ( .A1(n11466), .A2(n16387), .ZN(n7899) );
NOR2_X1 U25450 ( .A1(n10746), .A2(n16389), .ZN(n7869) );
NOR2_X1 U25451 ( .A1(n10745), .A2(n16387), .ZN(n7873) );
NOR2_X1 U25452 ( .A1(n10732), .A2(n16389), .ZN(n7879) );
NOR2_X1 U25453 ( .A1(n10731), .A2(n16387), .ZN(n7881) );
NOR2_X1 U25454 ( .A1(n10718), .A2(n16389), .ZN(n7891) );
NOR2_X1 U25455 ( .A1(n10717), .A2(n16387), .ZN(n7893) );
NOR2_X1 U25456 ( .A1(n10705), .A2(n16389), .ZN(n7903) );
NOR2_X1 U25457 ( .A1(n10704), .A2(n16387), .ZN(n7905) );
NOR2_X1 U25458 ( .A1(n10681), .A2(n16389), .ZN(n7885) );
NOR2_X1 U25459 ( .A1(n10680), .A2(n16387), .ZN(n7887) );
NOR2_X1 U25460 ( .A1(n10671), .A2(n16389), .ZN(n7909) );
NOR2_X1 U25461 ( .A1(n10670), .A2(n16387), .ZN(n7911) );
NAND2_X1 U25462 ( .A1(n11290), .A2(n15888), .ZN(n5550) );
NOR2_X1 U25463 ( .A1(n11006), .A2(n19969), .ZN(n15251) );
NOR2_X1 U25464 ( .A1(n11005), .A2(n19969), .ZN(n15250) );
NOR2_X1 U25465 ( .A1(n11004), .A2(n19969), .ZN(n15249) );
NOR2_X1 U25466 ( .A1(n11003), .A2(n19969), .ZN(n15248) );
NOR2_X1 U25467 ( .A1(n11002), .A2(n19969), .ZN(n15247) );
NOR2_X1 U25468 ( .A1(n11001), .A2(n19969), .ZN(n15246) );
NOR2_X1 U25469 ( .A1(n11000), .A2(n19969), .ZN(n15245) );
NOR2_X1 U25470 ( .A1(n10999), .A2(n19969), .ZN(n15244) );
NOR2_X1 U25471 ( .A1(n10998), .A2(n19969), .ZN(n15243) );
NOR2_X1 U25472 ( .A1(n10997), .A2(n19969), .ZN(n15242) );
NOR2_X1 U25473 ( .A1(n10996), .A2(n19969), .ZN(n15241) );
NOR2_X1 U25474 ( .A1(n10995), .A2(n19969), .ZN(n15240) );
NOR2_X1 U25475 ( .A1(n10994), .A2(n19969), .ZN(n15239) );
NOR2_X1 U25476 ( .A1(n10993), .A2(n19969), .ZN(n15238) );
NOR2_X1 U25477 ( .A1(n10992), .A2(n19969), .ZN(n15237) );
NOR2_X1 U25478 ( .A1(n10991), .A2(n19969), .ZN(n15236) );
NOR2_X1 U25479 ( .A1(n10990), .A2(n19969), .ZN(n15235) );
NOR2_X1 U25480 ( .A1(n10989), .A2(n19969), .ZN(n15234) );
NOR2_X1 U25481 ( .A1(n10988), .A2(n19969), .ZN(n15233) );
NOR2_X1 U25482 ( .A1(n10987), .A2(n19969), .ZN(n15232) );
NOR2_X1 U25483 ( .A1(n10986), .A2(n19969), .ZN(n15231) );
NOR2_X1 U25484 ( .A1(n10984), .A2(n19969), .ZN(n15229) );
NAND2_X1 U25485 ( .A1(n21407), .A2(n21406), .ZN(n21491) );
NAND2_X1 U25486 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_fifo_i_add_146_B_1_), .A2(crash_dump_o_66_), .ZN(n21406) );
NAND2_X1 U25487 ( .A1(n21446), .A2(crash_dump_o_66_), .ZN(n21407) );
NAND2_X1 U25488 ( .A1(n11064), .A2(n15818), .ZN(n1326) );
NAND2_X1 U25489 ( .A1(n10329), .A2(n8426), .ZN(n5237) );
NOR2_X1 U25490 ( .A1(n11519), .A2(n10330), .ZN(n10329) );
NAND2_X1 U25491 ( .A1(id_stage_i_controller_i_enter_debug_mode_prio_q), .A2(n5194), .ZN(n5152) );
NAND2_X1 U25492 ( .A1(n20915), .A2(n5196), .ZN(n5194) );
NAND2_X1 U25493 ( .A1(n10226), .A2(n10227), .ZN(n10104) );
NOR2_X1 U25494 ( .A1(n15910), .A2(n10231), .ZN(n10226) );
NOR2_X1 U25495 ( .A1(n15912), .A2(n10229), .ZN(n10227) );
NAND2_X1 U25496 ( .A1(n11317), .A2(n11322), .ZN(n10231) );
NOR2_X1 U25497 ( .A1(n10979), .A2(n16394), .ZN(n7555) );
NOR2_X1 U25498 ( .A1(n10831), .A2(n16393), .ZN(n7515) );
NOR2_X1 U25499 ( .A1(n10816), .A2(n16394), .ZN(n7523) );
NOR2_X1 U25500 ( .A1(n10802), .A2(n16393), .ZN(n7531) );
NOR2_X1 U25501 ( .A1(n10787), .A2(n16394), .ZN(n7539) );
NOR2_X1 U25502 ( .A1(n10768), .A2(n16393), .ZN(n7547) );
NOR2_X1 U25503 ( .A1(n10753), .A2(n16394), .ZN(n7566) );
NAND2_X1 U25504 ( .A1(n10409), .A2(n11502), .ZN(n10274) );
NOR2_X1 U25505 ( .A1(n10377), .A2(n1440), .ZN(n10409) );
NOR2_X1 U25506 ( .A1(n11018), .A2(n3776), .ZN(n3965) );
NOR2_X1 U25507 ( .A1(n10834), .A2(n3776), .ZN(n3909) );
NOR2_X1 U25508 ( .A1(n10881), .A2(n3776), .ZN(n3864) );
NOR2_X1 U25509 ( .A1(n10941), .A2(n3776), .ZN(n3808) );
NOR2_X1 U25510 ( .A1(n10971), .A2(n3776), .ZN(n3785) );
NOR2_X1 U25511 ( .A1(n10638), .A2(n3776), .ZN(n3769) );
NAND2_X1 U25512 ( .A1(n2830), .A2(n2831), .ZN(n2591) );
NOR2_X1 U25513 ( .A1(n2835), .A2(n2836), .ZN(n2830) );
NOR2_X1 U25514 ( .A1(n2832), .A2(n2833), .ZN(n2831) );
NOR2_X1 U25515 ( .A1(n11361), .A2(n16448), .ZN(n2835) );
NAND2_X1 U25516 ( .A1(n22109), .A2(n22108), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_N221) );
OR2_X1 U25517 ( .A1(n22107), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_4), .ZN(n22109) );
NAND2_X1 U25518 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_4), .A2(n22107), .ZN(n22108) );
NAND2_X1 U25519 ( .A1(n11299), .A2(n15823), .ZN(n4959) );
NOR2_X1 U25520 ( .A1(n11476), .A2(n7041), .ZN(n7038) );
NOR2_X1 U25521 ( .A1(n10969), .A2(n7323), .ZN(n7418) );
NOR2_X1 U25522 ( .A1(n10954), .A2(n7323), .ZN(n7426) );
NOR2_X1 U25523 ( .A1(n10939), .A2(n7323), .ZN(n7434) );
NOR2_X1 U25524 ( .A1(n10924), .A2(n7323), .ZN(n7442) );
NOR2_X1 U25525 ( .A1(n10909), .A2(n7323), .ZN(n7450) );
NOR2_X1 U25526 ( .A1(n10894), .A2(n7323), .ZN(n7458) );
NOR2_X1 U25527 ( .A1(n10879), .A2(n7323), .ZN(n7474) );
NOR2_X1 U25528 ( .A1(n10864), .A2(n7323), .ZN(n7490) );
NOR2_X1 U25529 ( .A1(n10847), .A2(n7323), .ZN(n7498) );
NOR2_X1 U25530 ( .A1(n10662), .A2(n16392), .ZN(n7394) );
NOR2_X1 U25531 ( .A1(n10647), .A2(n16392), .ZN(n7506) );
NOR2_X1 U25532 ( .A1(n11465), .A2(n7323), .ZN(n7482) );
NOR2_X1 U25533 ( .A1(n10632), .A2(n7323), .ZN(n7410) );
NOR2_X1 U25534 ( .A1(n10622), .A2(n16392), .ZN(n7402) );
NOR2_X1 U25535 ( .A1(n11495), .A2(n7323), .ZN(n7466) );
NOR2_X1 U25536 ( .A1(n11505), .A2(n16392), .ZN(n7386) );
NOR2_X1 U25537 ( .A1(n11512), .A2(n7872), .ZN(n7915) );
NOR2_X1 U25538 ( .A1(n11467), .A2(n7876), .ZN(n7917) );
NOR2_X1 U25539 ( .A1(n11506), .A2(n7872), .ZN(n7921) );
NOR2_X1 U25540 ( .A1(n11505), .A2(n7876), .ZN(n7923) );
NOR2_X1 U25541 ( .A1(n11496), .A2(n7872), .ZN(n7981) );
NOR2_X1 U25542 ( .A1(n11495), .A2(n7876), .ZN(n7983) );
NOR2_X1 U25543 ( .A1(n11485), .A2(n7872), .ZN(n7993) );
NOR2_X1 U25544 ( .A1(n11465), .A2(n7876), .ZN(n7995) );
NOR2_X1 U25545 ( .A1(n11455), .A2(n3130), .ZN(n3158) );
NOR2_X1 U25546 ( .A1(n11454), .A2(n3130), .ZN(n3162) );
NOR2_X1 U25547 ( .A1(n11453), .A2(n3130), .ZN(n3170) );
NOR2_X1 U25548 ( .A1(n11452), .A2(n3130), .ZN(n3174) );
NOR2_X1 U25549 ( .A1(n11451), .A2(n16435), .ZN(n3178) );
NOR2_X1 U25550 ( .A1(n11450), .A2(n3130), .ZN(n3182) );
NOR2_X1 U25551 ( .A1(n11449), .A2(n16435), .ZN(n3186) );
NOR2_X1 U25552 ( .A1(n11448), .A2(n3130), .ZN(n3190) );
NOR2_X1 U25553 ( .A1(n11447), .A2(n16435), .ZN(n3194) );
NOR2_X1 U25554 ( .A1(n11446), .A2(n3130), .ZN(n3198) );
NOR2_X1 U25555 ( .A1(n11445), .A2(n16435), .ZN(n3202) );
NOR2_X1 U25556 ( .A1(n11444), .A2(n3130), .ZN(n3206) );
NOR2_X1 U25557 ( .A1(n11443), .A2(n16435), .ZN(n3214) );
NOR2_X1 U25558 ( .A1(n11442), .A2(n3130), .ZN(n3218) );
NOR2_X1 U25559 ( .A1(n11441), .A2(n16435), .ZN(n3222) );
NOR2_X1 U25560 ( .A1(n11433), .A2(n3130), .ZN(n3127) );
NOR2_X1 U25561 ( .A1(n11432), .A2(n3130), .ZN(n3133) );
NOR2_X1 U25562 ( .A1(n11431), .A2(n3130), .ZN(n3138) );
NOR2_X1 U25563 ( .A1(n11430), .A2(n3130), .ZN(n3142) );
NOR2_X1 U25564 ( .A1(n11429), .A2(n16435), .ZN(n3146) );
NOR2_X1 U25565 ( .A1(n11428), .A2(n3130), .ZN(n3150) );
NOR2_X1 U25566 ( .A1(n11427), .A2(n16435), .ZN(n3154) );
NOR2_X1 U25567 ( .A1(n11426), .A2(n3130), .ZN(n3166) );
NOR2_X1 U25568 ( .A1(n11425), .A2(n3130), .ZN(n3210) );
NOR2_X1 U25569 ( .A1(n11422), .A2(n16433), .ZN(n3291) );
NOR2_X1 U25570 ( .A1(n11421), .A2(n16433), .ZN(n3295) );
NOR2_X1 U25571 ( .A1(n11420), .A2(n16433), .ZN(n3303) );
NOR2_X1 U25572 ( .A1(n11419), .A2(n16433), .ZN(n3307) );
NOR2_X1 U25573 ( .A1(n11418), .A2(n3263), .ZN(n3311) );
NOR2_X1 U25574 ( .A1(n11417), .A2(n3263), .ZN(n3315) );
NOR2_X1 U25575 ( .A1(n11416), .A2(n3263), .ZN(n3319) );
NOR2_X1 U25576 ( .A1(n11415), .A2(n16433), .ZN(n3323) );
NOR2_X1 U25577 ( .A1(n11414), .A2(n3263), .ZN(n3327) );
NOR2_X1 U25578 ( .A1(n11413), .A2(n16433), .ZN(n3331) );
NOR2_X1 U25579 ( .A1(n11412), .A2(n3263), .ZN(n3335) );
NOR2_X1 U25580 ( .A1(n11411), .A2(n16433), .ZN(n3339) );
NOR2_X1 U25581 ( .A1(n11410), .A2(n3263), .ZN(n3347) );
NOR2_X1 U25582 ( .A1(n11409), .A2(n16433), .ZN(n3351) );
NOR2_X1 U25583 ( .A1(n11408), .A2(n3263), .ZN(n3356) );
NOR2_X1 U25584 ( .A1(n11400), .A2(n16433), .ZN(n3260) );
NOR2_X1 U25585 ( .A1(n11399), .A2(n16433), .ZN(n3266) );
NOR2_X1 U25586 ( .A1(n11398), .A2(n16433), .ZN(n3270) );
NOR2_X1 U25587 ( .A1(n11397), .A2(n16433), .ZN(n3274) );
NOR2_X1 U25588 ( .A1(n11396), .A2(n16433), .ZN(n3278) );
NOR2_X1 U25589 ( .A1(n11395), .A2(n16433), .ZN(n3282) );
NOR2_X1 U25590 ( .A1(n11394), .A2(n16433), .ZN(n3286) );
NOR2_X1 U25591 ( .A1(n11393), .A2(n16433), .ZN(n3299) );
NOR2_X1 U25592 ( .A1(n11392), .A2(n16433), .ZN(n3343) );
NOR2_X1 U25593 ( .A1(n11308), .A2(n16389), .ZN(n8047) );
NOR2_X1 U25594 ( .A1(n11307), .A2(n16387), .ZN(n8049) );
NOR2_X1 U25595 ( .A1(n10970), .A2(n7872), .ZN(n7945) );
NOR2_X1 U25596 ( .A1(n10969), .A2(n7876), .ZN(n7947) );
NOR2_X1 U25597 ( .A1(n10955), .A2(n7872), .ZN(n7951) );
NOR2_X1 U25598 ( .A1(n10954), .A2(n7876), .ZN(n7953) );
NOR2_X1 U25599 ( .A1(n10940), .A2(n7872), .ZN(n7957) );
NOR2_X1 U25600 ( .A1(n10939), .A2(n7876), .ZN(n7959) );
NOR2_X1 U25601 ( .A1(n10925), .A2(n16389), .ZN(n7963) );
NOR2_X1 U25602 ( .A1(n10924), .A2(n16387), .ZN(n7965) );
NOR2_X1 U25603 ( .A1(n10910), .A2(n7872), .ZN(n7969) );
NOR2_X1 U25604 ( .A1(n10909), .A2(n7876), .ZN(n7971) );
NOR2_X1 U25605 ( .A1(n10865), .A2(n7872), .ZN(n7999) );
NOR2_X1 U25606 ( .A1(n10864), .A2(n7876), .ZN(n8001) );
NOR2_X1 U25607 ( .A1(n10848), .A2(n16389), .ZN(n8005) );
NOR2_X1 U25608 ( .A1(n10847), .A2(n16387), .ZN(n8007) );
NOR2_X1 U25609 ( .A1(n10833), .A2(n7872), .ZN(n8017) );
NOR2_X1 U25610 ( .A1(n10832), .A2(n7876), .ZN(n8019) );
NOR2_X1 U25611 ( .A1(n10818), .A2(n16389), .ZN(n8023) );
NOR2_X1 U25612 ( .A1(n10817), .A2(n16387), .ZN(n8025) );
NOR2_X1 U25613 ( .A1(n10663), .A2(n16389), .ZN(n7927) );
NOR2_X1 U25614 ( .A1(n10662), .A2(n16387), .ZN(n7929) );
NOR2_X1 U25615 ( .A1(n10648), .A2(n7872), .ZN(n8011) );
NOR2_X1 U25616 ( .A1(n10647), .A2(n7876), .ZN(n8013) );
NOR2_X1 U25617 ( .A1(n10633), .A2(n7872), .ZN(n7939) );
NOR2_X1 U25618 ( .A1(n10632), .A2(n7876), .ZN(n7941) );
NOR2_X1 U25619 ( .A1(n10623), .A2(n16389), .ZN(n7933) );
NOR2_X1 U25620 ( .A1(n10622), .A2(n16387), .ZN(n7935) );
NOR2_X1 U25621 ( .A1(n11194), .A2(n4291), .ZN(n4739) );
NOR2_X1 U25622 ( .A1(n11196), .A2(n4291), .ZN(n4700) );
NOR2_X1 U25623 ( .A1(n11197), .A2(n4291), .ZN(n4679) );
NOR2_X1 U25624 ( .A1(n11198), .A2(n4291), .ZN(n4658) );
NOR2_X1 U25625 ( .A1(n11199), .A2(n4291), .ZN(n4637) );
NOR2_X1 U25626 ( .A1(n11200), .A2(n4291), .ZN(n4616) );
NOR2_X1 U25627 ( .A1(n11201), .A2(n4291), .ZN(n4595) );
NOR2_X1 U25628 ( .A1(n11202), .A2(n16419), .ZN(n4574) );
NOR2_X1 U25629 ( .A1(n11203), .A2(n4291), .ZN(n4553) );
NOR2_X1 U25630 ( .A1(n11204), .A2(n16419), .ZN(n4532) );
NOR2_X1 U25631 ( .A1(n11195), .A2(n4291), .ZN(n4719) );
NOR2_X1 U25632 ( .A1(n11214), .A2(n16419), .ZN(n4276) );
NOR2_X1 U25633 ( .A1(n11014), .A2(n6719), .ZN(n6813) );
NOR2_X1 U25634 ( .A1(n11012), .A2(n16402), .ZN(n6915) );
NOR2_X1 U25635 ( .A1(n11011), .A2(n16402), .ZN(n6991) );
NOR2_X1 U25636 ( .A1(n11010), .A2(n16402), .ZN(n7001) );
NOR2_X1 U25637 ( .A1(n11009), .A2(n6719), .ZN(n7026) );
NOR2_X1 U25638 ( .A1(n10895), .A2(n7872), .ZN(n7975) );
NOR2_X1 U25639 ( .A1(n10894), .A2(n7876), .ZN(n7977) );
NOR2_X1 U25640 ( .A1(n10880), .A2(n16389), .ZN(n7987) );
NOR2_X1 U25641 ( .A1(n10879), .A2(n16387), .ZN(n7989) );
NOR2_X1 U25642 ( .A1(n10821), .A2(n16402), .ZN(n6961) );
NOR2_X1 U25643 ( .A1(n10804), .A2(n7872), .ZN(n8029) );
NOR2_X1 U25644 ( .A1(n10803), .A2(n7876), .ZN(n8031) );
NOR2_X1 U25645 ( .A1(n10788), .A2(n16387), .ZN(n8037) );
NOR2_X1 U25646 ( .A1(n10806), .A2(n16402), .ZN(n6971) );
NOR2_X1 U25647 ( .A1(n10789), .A2(n16389), .ZN(n8035) );
NOR2_X1 U25648 ( .A1(n10792), .A2(n16402), .ZN(n6981) );
NOR2_X1 U25649 ( .A1(n10770), .A2(n7872), .ZN(n8041) );
NOR2_X1 U25650 ( .A1(n10769), .A2(n7876), .ZN(n8043) );
NOR2_X1 U25651 ( .A1(n10760), .A2(n16389), .ZN(n8053) );
NOR2_X1 U25652 ( .A1(n10759), .A2(n16387), .ZN(n8057) );
NOR2_X1 U25653 ( .A1(n10754), .A2(n16402), .ZN(n7011) );
NOR2_X1 U25654 ( .A1(n10740), .A2(n16402), .ZN(n6713) );
NOR2_X1 U25655 ( .A1(n11332), .A2(n16451), .ZN(n2154) );
NOR2_X1 U25656 ( .A1(n11304), .A2(n20924), .ZN(n7063) );
NOR2_X1 U25657 ( .A1(n10778), .A2(n16354), .ZN(n7055) );
NOR2_X1 U25658 ( .A1(n10738), .A2(n20924), .ZN(n7314) );
NOR2_X1 U25659 ( .A1(n11217), .A2(n4291), .ZN(n4920) );
NOR2_X1 U25660 ( .A1(n11215), .A2(n16419), .ZN(n4450) );
NOR2_X1 U25661 ( .A1(n11205), .A2(n4291), .ZN(n4511) );
NOR2_X1 U25662 ( .A1(n11207), .A2(n16419), .ZN(n4471) );
NOR2_X1 U25663 ( .A1(n11206), .A2(n4291), .ZN(n4490) );
NOR2_X1 U25664 ( .A1(n11208), .A2(n16419), .ZN(n4396) );
NOR2_X1 U25665 ( .A1(n11209), .A2(n4291), .ZN(n4377) );
NOR2_X1 U25666 ( .A1(n11210), .A2(n16419), .ZN(n4358) );
NOR2_X1 U25667 ( .A1(n11211), .A2(n4291), .ZN(n4339) );
NOR2_X1 U25668 ( .A1(n11212), .A2(n16419), .ZN(n4320) );
NOR2_X1 U25669 ( .A1(n11213), .A2(n4291), .ZN(n4301) );
NAND2_X1 U25670 ( .A1(n5227), .A2(n5228), .ZN(n5178) );
NOR2_X1 U25671 ( .A1(n15800), .A2(n15915), .ZN(n5227) );
NOR2_X1 U25672 ( .A1(n11514), .A2(n15798), .ZN(n5228) );
NOR2_X1 U25673 ( .A1(n11305), .A2(n7041), .ZN(n8139) );
NOR2_X1 U25674 ( .A1(n10779), .A2(n7041), .ZN(n8134) );
NOR2_X1 U25675 ( .A1(n19814), .A2(n6552), .ZN(n6565) );
INV_X1 U25676 ( .A(boot_addr_i_31_), .ZN(n19814) );
NOR2_X1 U25677 ( .A1(n19816), .A2(n6552), .ZN(n6571) );
INV_X1 U25678 ( .A(boot_addr_i_30_), .ZN(n19816) );
NOR2_X1 U25679 ( .A1(n19819), .A2(n16404), .ZN(n6577) );
INV_X1 U25680 ( .A(boot_addr_i_29_), .ZN(n19819) );
NOR2_X1 U25681 ( .A1(n19839), .A2(n6552), .ZN(n6625) );
INV_X1 U25682 ( .A(boot_addr_i_21_), .ZN(n19839) );
NOR2_X1 U25683 ( .A1(n19864), .A2(n16404), .ZN(n6685) );
INV_X1 U25684 ( .A(boot_addr_i_11_), .ZN(n19864) );
NOR2_X1 U25685 ( .A1(n19824), .A2(n6552), .ZN(n6589) );
INV_X1 U25686 ( .A(boot_addr_i_27_), .ZN(n19824) );
NOR2_X1 U25687 ( .A1(n19827), .A2(n16404), .ZN(n6595) );
INV_X1 U25688 ( .A(boot_addr_i_26_), .ZN(n19827) );
NOR2_X1 U25689 ( .A1(n19829), .A2(n6552), .ZN(n6601) );
INV_X1 U25690 ( .A(boot_addr_i_25_), .ZN(n19829) );
NOR2_X1 U25691 ( .A1(n19832), .A2(n16404), .ZN(n6607) );
INV_X1 U25692 ( .A(boot_addr_i_24_), .ZN(n19832) );
NOR2_X1 U25693 ( .A1(n19834), .A2(n6552), .ZN(n6613) );
INV_X1 U25694 ( .A(boot_addr_i_23_), .ZN(n19834) );
NOR2_X1 U25695 ( .A1(n19837), .A2(n16404), .ZN(n6619) );
INV_X1 U25696 ( .A(boot_addr_i_22_), .ZN(n19837) );
NOR2_X1 U25697 ( .A1(n19842), .A2(n6552), .ZN(n6631) );
INV_X1 U25698 ( .A(boot_addr_i_20_), .ZN(n19842) );
NOR2_X1 U25699 ( .A1(n19844), .A2(n16404), .ZN(n6637) );
INV_X1 U25700 ( .A(boot_addr_i_19_), .ZN(n19844) );
NOR2_X1 U25701 ( .A1(n19847), .A2(n6552), .ZN(n6643) );
INV_X1 U25702 ( .A(boot_addr_i_18_), .ZN(n19847) );
NOR2_X1 U25703 ( .A1(n19852), .A2(n16404), .ZN(n6655) );
INV_X1 U25704 ( .A(boot_addr_i_16_), .ZN(n19852) );
NOR2_X1 U25705 ( .A1(n19854), .A2(n6552), .ZN(n6661) );
INV_X1 U25706 ( .A(boot_addr_i_15_), .ZN(n19854) );
NOR2_X1 U25707 ( .A1(n19857), .A2(n16404), .ZN(n6667) );
INV_X1 U25708 ( .A(boot_addr_i_14_), .ZN(n19857) );
NOR2_X1 U25709 ( .A1(n19859), .A2(n6552), .ZN(n6673) );
INV_X1 U25710 ( .A(boot_addr_i_13_), .ZN(n19859) );
NOR2_X1 U25711 ( .A1(n19862), .A2(n16404), .ZN(n6679) );
INV_X1 U25712 ( .A(boot_addr_i_12_), .ZN(n19862) );
NOR2_X1 U25713 ( .A1(n19867), .A2(n6552), .ZN(n6691) );
INV_X1 U25714 ( .A(boot_addr_i_10_), .ZN(n19867) );
NOR2_X1 U25715 ( .A1(n19869), .A2(n6552), .ZN(n6550) );
INV_X1 U25716 ( .A(boot_addr_i_9_), .ZN(n19869) );
NOR2_X1 U25717 ( .A1(n19872), .A2(n16404), .ZN(n6558) );
INV_X1 U25718 ( .A(boot_addr_i_8_), .ZN(n19872) );
NOR2_X1 U25719 ( .A1(n19849), .A2(n16404), .ZN(n6649) );
INV_X1 U25720 ( .A(boot_addr_i_17_), .ZN(n19849) );
NOR2_X1 U25721 ( .A1(n19822), .A2(n6552), .ZN(n6583) );
INV_X1 U25722 ( .A(boot_addr_i_28_), .ZN(n19822) );
NOR2_X1 U25723 ( .A1(n11330), .A2(n16452), .ZN(n2240) );
NAND2_X1 U25724 ( .A1(n11289), .A2(n15888), .ZN(n4926) );
NOR2_X1 U25725 ( .A1(n11379), .A2(n2169), .ZN(n2230) );
NOR2_X1 U25726 ( .A1(n2547), .A2(n2548), .ZN(n2546) );
NAND2_X1 U25727 ( .A1(n2549), .A2(n2550), .ZN(n2548) );
NOR2_X1 U25728 ( .A1(n11387), .A2(n16448), .ZN(n2547) );
NAND2_X1 U25729 ( .A1(instr_rdata_i_29_), .A2(n16447), .ZN(n2549) );
NAND2_X1 U25730 ( .A1(n1579), .A2(n16145), .ZN(n1550) );
NOR2_X1 U25731 ( .A1(n11469), .A2(n19886), .ZN(n3719) );
NOR2_X1 U25732 ( .A1(n11424), .A2(n3263), .ZN(n3390) );
NOR2_X1 U25733 ( .A1(n11407), .A2(n3263), .ZN(n3361) );
NOR2_X1 U25734 ( .A1(n11406), .A2(n3263), .ZN(n3365) );
NOR2_X1 U25735 ( .A1(n11405), .A2(n3263), .ZN(n3369) );
NOR2_X1 U25736 ( .A1(n11404), .A2(n3263), .ZN(n3373) );
NOR2_X1 U25737 ( .A1(n11403), .A2(n3263), .ZN(n3377) );
NOR2_X1 U25738 ( .A1(n11402), .A2(n3263), .ZN(n3381) );
NOR2_X1 U25739 ( .A1(n11401), .A2(n3263), .ZN(n3385) );
NOR2_X1 U25740 ( .A1(n11457), .A2(n16435), .ZN(n3255) );
NOR2_X1 U25741 ( .A1(n11440), .A2(n16435), .ZN(n3227) );
NOR2_X1 U25742 ( .A1(n11439), .A2(n16435), .ZN(n3231) );
NOR2_X1 U25743 ( .A1(n11438), .A2(n16435), .ZN(n3235) );
NOR2_X1 U25744 ( .A1(n11437), .A2(n16435), .ZN(n3239) );
NOR2_X1 U25745 ( .A1(n11436), .A2(n16435), .ZN(n3243) );
NOR2_X1 U25746 ( .A1(n11435), .A2(n16435), .ZN(n3247) );
NOR2_X1 U25747 ( .A1(n11434), .A2(n16435), .ZN(n3251) );
NOR2_X1 U25748 ( .A1(n11016), .A2(n6719), .ZN(n6759) );
NOR2_X1 U25749 ( .A1(n11015), .A2(n6719), .ZN(n6781) );
NOR2_X1 U25750 ( .A1(n10726), .A2(n6719), .ZN(n6726) );
NOR2_X1 U25751 ( .A1(n10712), .A2(n6719), .ZN(n6748) );
NOR2_X1 U25752 ( .A1(n10699), .A2(n6719), .ZN(n6770) );
NOR2_X1 U25753 ( .A1(n10687), .A2(n6719), .ZN(n6737) );
NOR2_X1 U25754 ( .A1(n2736), .A2(n2737), .ZN(n2735) );
NOR2_X1 U25755 ( .A1(n15803), .A2(n2738), .ZN(n2736) );
NOR2_X1 U25756 ( .A1(n11423), .A2(n2164), .ZN(n2737) );
NAND2_X1 U25757 ( .A1(n20903), .A2(n19962), .ZN(n2738) );
NOR2_X1 U25758 ( .A1(n1554), .A2(n1699), .ZN(n1693) );
NAND2_X1 U25759 ( .A1(data_rvalid_i), .A2(n20022), .ZN(n1699) );
NOR2_X1 U25760 ( .A1(n11329), .A2(n15858), .ZN(n10395) );
NOR2_X1 U25761 ( .A1(n5245), .A2(n5246), .ZN(n5243) );
NOR2_X1 U25762 ( .A1(n5247), .A2(n5248), .ZN(n5246) );
NOR2_X1 U25763 ( .A1(n5249), .A2(n5250), .ZN(n5248) );
NOR2_X1 U25764 ( .A1(n11499), .A2(n5173), .ZN(n5247) );
NOR2_X1 U25765 ( .A1(n1571), .A2(n1692), .ZN(n1691) );
NAND2_X1 U25766 ( .A1(n11294), .A2(n1549), .ZN(n1692) );
NOR2_X1 U25767 ( .A1(n4432), .A2(n4433), .ZN(n4430) );
NOR2_X1 U25768 ( .A1(n11216), .A2(n4435), .ZN(n4432) );
NOR2_X1 U25769 ( .A1(n20110), .A2(n20112), .ZN(n4433) );
NOR2_X1 U25770 ( .A1(n10250), .A2(n10251), .ZN(n10249) );
NAND2_X1 U25771 ( .A1(n10252), .A2(n11333), .ZN(n10251) );
NAND2_X1 U25772 ( .A1(n10254), .A2(n10255), .ZN(n10250) );
NOR2_X1 U25773 ( .A1(n10253), .A2(n15860), .ZN(n10252) );
NOR2_X1 U25774 ( .A1(n3056), .A2(n3018), .ZN(n3052) );
NOR2_X1 U25775 ( .A1(n3057), .A2(n3058), .ZN(n3056) );
NOR2_X1 U25776 ( .A1(n11459), .A2(n19884), .ZN(n3057) );
NOR2_X1 U25777 ( .A1(n11460), .A2(n3042), .ZN(n3058) );
NOR2_X1 U25778 ( .A1(n11320), .A2(n1596), .ZN(n10407) );
NOR2_X1 U25779 ( .A1(n11312), .A2(n15859), .ZN(n10261) );
NOR2_X1 U25780 ( .A1(n11500), .A2(n5113), .ZN(n5109) );
NOR2_X1 U25781 ( .A1(n19987), .A2(n1431), .ZN(n5113) );
INV_X1 U25782 ( .A(n5115), .ZN(n19987) );
NOR2_X1 U25783 ( .A1(n11298), .A2(n1531), .ZN(n1551) );
NOR2_X1 U25784 ( .A1(n11477), .A2(n16399), .ZN(n7044) );
NOR2_X1 U25785 ( .A1(n11459), .A2(n16116), .ZN(n2660) );
NOR2_X1 U25786 ( .A1(n11459), .A2(n16117), .ZN(n2503) );
NOR2_X1 U25787 ( .A1(n11459), .A2(n16118), .ZN(n2296) );
NAND2_X1 U25788 ( .A1(n10297), .A2(n11314), .ZN(n10253) );
NOR2_X1 U25789 ( .A1(n15827), .A2(n16119), .ZN(n10297) );
NOR2_X1 U25790 ( .A1(n1540), .A2(n1541), .ZN(n1539) );
NOR2_X1 U25791 ( .A1(n1542), .A2(n1543), .ZN(n1540) );
AND2_X1 U25792 ( .A1(n1544), .A2(data_gnt_i), .ZN(n1542) );
NOR2_X1 U25793 ( .A1(data_gnt_i), .A2(n1544), .ZN(n1543) );
NOR2_X1 U25794 ( .A1(n10078), .A2(n10079), .ZN(n10077) );
OR2_X1 U25795 ( .A1(n6509), .A2(n11519), .ZN(n10079) );
NOR2_X1 U25796 ( .A1(n1575), .A2(n10080), .ZN(n10078) );
NAND2_X1 U25797 ( .A1(n1444), .A2(n1580), .ZN(n10080) );
NOR2_X1 U25798 ( .A1(n10381), .A2(n10382), .ZN(n10380) );
NAND2_X1 U25799 ( .A1(n10383), .A2(n15804), .ZN(n10382) );
NOR2_X1 U25800 ( .A1(n11501), .A2(n11502), .ZN(n10381) );
NAND2_X1 U25801 ( .A1(n10384), .A2(n10385), .ZN(n10383) );
NOR2_X1 U25802 ( .A1(n11321), .A2(n15908), .ZN(n10534) );
NOR2_X1 U25803 ( .A1(n11165), .A2(n4946), .ZN(n4945) );
NOR2_X1 U25804 ( .A1(n20910), .A2(n4947), .ZN(n4946) );
NAND2_X1 U25805 ( .A1(n4797), .A2(n4918), .ZN(n4947) );
AND2_X1 U25806 ( .A1(n5263), .A2(n10434), .ZN(n8426) );
NOR2_X1 U25807 ( .A1(rf_raddr_b_o_2_), .A2(n10435), .ZN(n10434) );
NAND2_X1 U25808 ( .A1(n11338), .A2(n10287), .ZN(n10435) );
AND2_X1 U25809 ( .A1(n5097), .A2(n5098), .ZN(n4423) );
NAND2_X1 U25810 ( .A1(n5099), .A2(n11219), .ZN(n5098) );
NAND2_X1 U25811 ( .A1(n20085), .A2(n4940), .ZN(n5097) );
NOR2_X1 U25812 ( .A1(n5100), .A2(n4940), .ZN(n5099) );
NAND2_X1 U25813 ( .A1(n11293), .A2(n6532), .ZN(n6525) );
OR2_X1 U25814 ( .A1(n1565), .A2(n1590), .ZN(n6532) );
OR2_X1 U25815 ( .A1(n16272), .A2(n1440), .ZN(n1439) );
OR2_X1 U25816 ( .A1(n11502), .A2(n10377), .ZN(n16272) );
AND2_X1 U25817 ( .A1(n10327), .A2(n10548), .ZN(n7712) );
NOR2_X1 U25818 ( .A1(n5238), .A2(n10328), .ZN(n10327) );
NOR2_X1 U25819 ( .A1(rf_raddr_b_o_0_), .A2(n5237), .ZN(n10328) );
NOR2_X1 U25820 ( .A1(n2226), .A2(n2227), .ZN(n2225) );
NOR2_X1 U25821 ( .A1(n19957), .A2(n2166), .ZN(n2226) );
NOR2_X1 U25822 ( .A1(n11395), .A2(n2164), .ZN(n2227) );
NAND2_X1 U25823 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_31), .ZN(n4452) );
NAND2_X1 U25824 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_3), .ZN(n4398) );
NAND2_X1 U25825 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_4), .ZN(n4379) );
NAND2_X1 U25826 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_5), .ZN(n4360) );
NAND2_X1 U25827 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_6), .ZN(n4341) );
NAND2_X1 U25828 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_7), .ZN(n4322) );
NAND2_X1 U25829 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_8), .ZN(n4303) );
NOR2_X1 U25830 ( .A1(n11320), .A2(n15895), .ZN(n10385) );
NAND2_X1 U25831 ( .A1(n10324), .A2(n10325), .ZN(n5196) );
NAND2_X1 U25832 ( .A1(n10326), .A2(n16042), .ZN(n10325) );
NAND2_X1 U25833 ( .A1(n5245), .A2(n16043), .ZN(n10324) );
NOR2_X1 U25834 ( .A1(priv_mode_id_1), .A2(priv_mode_id_0), .ZN(n10326) );
NAND2_X1 U25835 ( .A1(crash_dump_o_125_), .A2(n20899), .ZN(n21594) );
INV_X1 U25836 ( .A(n21591), .ZN(n20899) );
NAND2_X1 U25837 ( .A1(crash_dump_o_93_), .A2(n19937), .ZN(n21487) );
INV_X1 U25838 ( .A(n21482), .ZN(n19937) );
NAND2_X1 U25839 ( .A1(cs_registers_i_mhpmcounter_2__61_), .A2(n20901), .ZN(n22529) );
INV_X1 U25840 ( .A(n22526), .ZN(n20901) );
NAND2_X1 U25841 ( .A1(cs_registers_i_mhpmcounter_0__61_), .A2(n20897), .ZN(n22311) );
INV_X1 U25842 ( .A(n22308), .ZN(n20897) );
NAND2_X1 U25843 ( .A1(n21585), .A2(crash_dump_o_124_), .ZN(n21591) );
NOR2_X1 U25844 ( .A1(n21584), .A2(n10969), .ZN(n21585) );
NAND2_X1 U25845 ( .A1(n21479), .A2(crash_dump_o_92_), .ZN(n21482) );
NOR2_X1 U25846 ( .A1(n21478), .A2(n10970), .ZN(n21479) );
NAND2_X1 U25847 ( .A1(n22523), .A2(cs_registers_i_mhpmcounter_2__60_), .ZN(n22526) );
NOR2_X1 U25848 ( .A1(n22522), .A2(n10966), .ZN(n22523) );
NAND2_X1 U25849 ( .A1(n22305), .A2(cs_registers_i_mhpmcounter_0__60_), .ZN(n22308) );
NOR2_X1 U25850 ( .A1(n22304), .A2(n10964), .ZN(n22305) );
NAND2_X1 U25851 ( .A1(n10466), .A2(n10461), .ZN(n5168) );
NOR2_X1 U25852 ( .A1(n11517), .A2(n15798), .ZN(n10466) );
NAND2_X1 U25853 ( .A1(n3718), .A2(n15929), .ZN(n3710) );
NAND2_X1 U25854 ( .A1(n11470), .A2(n16439), .ZN(n3718) );
NOR2_X1 U25855 ( .A1(n7663), .A2(n7664), .ZN(n7636) );
NOR2_X1 U25856 ( .A1(n19809), .A2(n7562), .ZN(n7663) );
NOR2_X1 U25857 ( .A1(n11487), .A2(n16354), .ZN(n7664) );
NOR2_X1 U25858 ( .A1(n7631), .A2(n7632), .ZN(n7611) );
NOR2_X1 U25859 ( .A1(n19807), .A2(n7562), .ZN(n7631) );
NOR2_X1 U25860 ( .A1(n11481), .A2(n16354), .ZN(n7632) );
NOR2_X1 U25861 ( .A1(n7714), .A2(n7715), .ZN(n7668) );
NOR2_X1 U25862 ( .A1(n19811), .A2(n7562), .ZN(n7714) );
NOR2_X1 U25863 ( .A1(n10854), .A2(n16354), .ZN(n7715) );
NOR2_X1 U25864 ( .A1(n7606), .A2(n7607), .ZN(n7595) );
NOR2_X1 U25865 ( .A1(n19805), .A2(n7562), .ZN(n7606) );
NOR2_X1 U25866 ( .A1(n10676), .A2(n16354), .ZN(n7607) );
NAND2_X1 U25867 ( .A1(n11299), .A2(n11300), .ZN(n5087) );
NOR2_X1 U25868 ( .A1(n10404), .A2(n10405), .ZN(n10399) );
NOR2_X1 U25869 ( .A1(n11329), .A2(n10406), .ZN(n10405) );
NOR2_X1 U25870 ( .A1(n10412), .A2(n10070), .ZN(n10404) );
NOR2_X1 U25871 ( .A1(n10407), .A2(n20976), .ZN(n10406) );
NOR2_X1 U25872 ( .A1(n10488), .A2(n10489), .ZN(n10486) );
AND2_X1 U25873 ( .A1(n10481), .A2(rf_waddr_wb_o_2_), .ZN(n10489) );
NOR2_X1 U25874 ( .A1(n20966), .A2(n10491), .ZN(n10488) );
NOR2_X1 U25875 ( .A1(n10492), .A2(n10156), .ZN(n10491) );
NOR2_X1 U25876 ( .A1(n2747), .A2(n2748), .ZN(n2744) );
NOR2_X1 U25877 ( .A1(n11390), .A2(n2754), .ZN(n2747) );
NOR2_X1 U25878 ( .A1(n2749), .A2(n2750), .ZN(n2748) );
NOR2_X1 U25879 ( .A1(n20903), .A2(n2755), .ZN(n2754) );
NOR2_X1 U25880 ( .A1(n10054), .A2(n10055), .ZN(n10052) );
NOR2_X1 U25881 ( .A1(n11316), .A2(n10056), .ZN(n10055) );
NOR2_X1 U25882 ( .A1(n16123), .A2(n10060), .ZN(n10054) );
NOR2_X1 U25883 ( .A1(n20954), .A2(n20955), .ZN(n10056) );
NOR2_X1 U25884 ( .A1(n10258), .A2(n10259), .ZN(n10254) );
NOR2_X1 U25885 ( .A1(n11339), .A2(n10260), .ZN(n10259) );
NOR2_X1 U25886 ( .A1(n10097), .A2(n10262), .ZN(n10258) );
NOR2_X1 U25887 ( .A1(n10261), .A2(n15816), .ZN(n10260) );
NOR2_X1 U25888 ( .A1(n11321), .A2(n15814), .ZN(n10242) );
INV_X1 U25889 ( .A(instr_rdata_i_30_), .ZN(n19911) );
INV_X1 U25890 ( .A(instr_rdata_i_29_), .ZN(n19913) );
INV_X1 U25891 ( .A(instr_rdata_i_25_), .ZN(n19922) );
INV_X1 U25892 ( .A(instr_rdata_i_24_), .ZN(n19924) );
INV_X1 U25893 ( .A(instr_rdata_i_22_), .ZN(n19928) );
INV_X1 U25894 ( .A(instr_rdata_i_21_), .ZN(n19930) );
INV_X1 U25895 ( .A(instr_rdata_i_19_), .ZN(n19933) );
INV_X1 U25896 ( .A(instr_rdata_i_14_), .ZN(n19947) );
INV_X1 U25897 ( .A(instr_rdata_i_13_), .ZN(n19948) );
INV_X1 U25898 ( .A(instr_rdata_i_8_), .ZN(n19953) );
INV_X1 U25899 ( .A(instr_rdata_i_6_), .ZN(n19955) );
INV_X1 U25900 ( .A(instr_rdata_i_5_), .ZN(n19956) );
INV_X1 U25901 ( .A(instr_rdata_i_3_), .ZN(n19958) );
NOR2_X1 U25902 ( .A1(n11313), .A2(n10369), .ZN(n10368) );
NOR2_X1 U25903 ( .A1(n10370), .A2(n10286), .ZN(n10369) );
NAND2_X1 U25904 ( .A1(n10287), .A2(n11325), .ZN(n10370) );
NOR2_X1 U25905 ( .A1(n11291), .A2(n5035), .ZN(n4978) );
NOR2_X1 U25906 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N221), .A2(n5036), .ZN(n5035) );
NOR2_X1 U25907 ( .A1(n5037), .A2(n5038), .ZN(n5036) );
NOR2_X1 U25908 ( .A1(n5039), .A2(n21011), .ZN(n5038) );
NOR2_X1 U25909 ( .A1(n11313), .A2(n11340), .ZN(n10366) );
NOR2_X1 U25910 ( .A1(n11338), .A2(n11493), .ZN(n5259) );
NAND2_X1 U25911 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_11), .ZN(n4900) );
NAND2_X1 U25912 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_12), .ZN(n4881) );
NAND2_X1 U25913 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_13), .ZN(n4862) );
NAND2_X1 U25914 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_14), .ZN(n4843) );
NAND2_X1 U25915 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_15), .ZN(n4824) );
NAND2_X1 U25916 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_16), .ZN(n4805) );
NAND2_X1 U25917 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_17), .ZN(n4783) );
NAND2_X1 U25918 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_18), .ZN(n4762) );
NAND2_X1 U25919 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_19), .ZN(n4741) );
NAND2_X1 U25920 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_1), .ZN(n4721) );
NAND2_X1 U25921 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_9), .ZN(n4278) );
NAND2_X1 U25922 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_10), .ZN(n4922) );
NAND2_X1 U25923 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_20), .ZN(n4702) );
NAND2_X1 U25924 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_21), .ZN(n4681) );
NAND2_X1 U25925 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_22), .ZN(n4660) );
NAND2_X1 U25926 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_23), .ZN(n4639) );
NAND2_X1 U25927 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_24), .ZN(n4618) );
NAND2_X1 U25928 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_25), .ZN(n4597) );
NAND2_X1 U25929 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_26), .ZN(n4576) );
NAND2_X1 U25930 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_27), .ZN(n4555) );
NAND2_X1 U25931 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_28), .ZN(n4534) );
NAND2_X1 U25932 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_29), .ZN(n4513) );
NAND2_X1 U25933 ( .A1(n20909), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_30), .ZN(n4473) );
NAND2_X1 U25934 ( .A1(n16352), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_2), .ZN(n4492) );
NAND2_X1 U25935 ( .A1(n11291), .A2(n4940), .ZN(n4932) );
OR2_X1 U25936 ( .A1(n10548), .A2(n5238), .ZN(n7025) );
NAND2_X1 U25937 ( .A1(n11485), .A2(n15793), .ZN(n2169) );
AND2_X1 U25938 ( .A1(n10067), .A2(n20937), .ZN(n9958) );
NOR2_X1 U25939 ( .A1(n11313), .A2(n10066), .ZN(n10067) );
NAND2_X1 U25940 ( .A1(n11485), .A2(n11460), .ZN(n2170) );
NAND2_X1 U25941 ( .A1(n16388), .A2(crash_dump_o_96_), .ZN(n8063) );
NAND2_X1 U25942 ( .A1(n10531), .A2(n10230), .ZN(n10248) );
NOR2_X1 U25943 ( .A1(n10532), .A2(n10533), .ZN(n10531) );
NOR2_X1 U25944 ( .A1(n11321), .A2(n10150), .ZN(n10533) );
NOR2_X1 U25945 ( .A1(n11317), .A2(n10534), .ZN(n10532) );
NAND2_X1 U25946 ( .A1(n10236), .A2(n10237), .ZN(n10148) );
NOR2_X1 U25947 ( .A1(n10247), .A2(n10248), .ZN(n10236) );
NOR2_X1 U25948 ( .A1(n10238), .A2(n10239), .ZN(n10237) );
NOR2_X1 U25949 ( .A1(n11322), .A2(n15910), .ZN(n10247) );
NAND2_X1 U25950 ( .A1(n11297), .A2(n20022), .ZN(n1698) );
NAND2_X1 U25951 ( .A1(n10454), .A2(n10455), .ZN(n10438) );
NOR2_X1 U25952 ( .A1(n11493), .A2(rf_raddr_b_o_0_), .ZN(n10454) );
NOR2_X1 U25953 ( .A1(n11331), .A2(n11338), .ZN(n10455) );
OR2_X1 U25954 ( .A1(n16273), .A2(n5141), .ZN(n5130) );
NAND2_X1 U25955 ( .A1(n5142), .A2(n11515), .ZN(n16273) );
NAND2_X1 U25956 ( .A1(n10522), .A2(n11327), .ZN(n10246) );
NOR2_X1 U25957 ( .A1(n11317), .A2(n10523), .ZN(n10522) );
NAND2_X1 U25958 ( .A1(n10530), .A2(n11321), .ZN(n9968) );
NOR2_X1 U25959 ( .A1(n11327), .A2(n10248), .ZN(n10530) );
NAND2_X1 U25960 ( .A1(n7707), .A2(n7708), .ZN(n7605) );
AND2_X1 U25961 ( .A1(n20923), .A2(n10548), .ZN(n7707) );
NOR2_X1 U25962 ( .A1(n5238), .A2(rf_raddr_b_o_0_), .ZN(n7708) );
NAND2_X1 U25963 ( .A1(n7662), .A2(n7710), .ZN(n7630) );
NAND2_X1 U25964 ( .A1(n7711), .A2(n7712), .ZN(n7710) );
NOR2_X1 U25965 ( .A1(n10547), .A2(n20923), .ZN(n7711) );
NAND2_X1 U25966 ( .A1(n4926), .A2(n6228), .ZN(n6222) );
NAND2_X1 U25967 ( .A1(n11290), .A2(n15887), .ZN(n6228) );
NAND2_X1 U25968 ( .A1(n10257), .A2(n11324), .ZN(n10187) );
NOR2_X1 U25969 ( .A1(n15860), .A2(n5580), .ZN(n10257) );
NAND2_X1 U25970 ( .A1(n5559), .A2(n5560), .ZN(n5542) );
AND2_X1 U25971 ( .A1(n11253), .A2(n11252), .ZN(n5559) );
NOR2_X1 U25972 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_2), .A2(n5562), .ZN(n5560) );
NAND2_X1 U25973 ( .A1(n10538), .A2(n11298), .ZN(n1581) );
NOR2_X1 U25974 ( .A1(n11296), .A2(n15925), .ZN(n10538) );
NAND2_X1 U25975 ( .A1(n11064), .A2(n1326), .ZN(n1359) );
NAND2_X1 U25976 ( .A1(n10278), .A2(n10279), .ZN(n10272) );
NOR2_X1 U25977 ( .A1(n5736), .A2(n20992), .ZN(n10279) );
NOR2_X1 U25978 ( .A1(n16357), .A2(n10291), .ZN(n10278) );
AND2_X1 U25979 ( .A1(n4426), .A2(n11291), .ZN(n10291) );
NOR2_X1 U25980 ( .A1(n11464), .A2(n8773), .ZN(n9962) );
NAND2_X1 U25981 ( .A1(n3597), .A2(n3598), .ZN(n2863) );
NAND2_X1 U25982 ( .A1(instr_rdata_i_17_), .A2(n11460), .ZN(n3598) );
NAND2_X1 U25983 ( .A1(n15793), .A2(n16044), .ZN(n3597) );
NAND2_X1 U25984 ( .A1(n2656), .A2(n2657), .ZN(n2644) );
NAND2_X1 U25985 ( .A1(instr_rdata_i_25_), .A2(n16447), .ZN(n2657) );
NOR2_X1 U25986 ( .A1(n2658), .A2(n2659), .ZN(n2656) );
NOR2_X1 U25987 ( .A1(n2660), .A2(n2661), .ZN(n2658) );
NAND2_X1 U25988 ( .A1(n2662), .A2(crash_dump_o_65_), .ZN(n2661) );
NAND2_X1 U25989 ( .A1(n11459), .A2(n19952), .ZN(n2662) );
NAND2_X1 U25990 ( .A1(n2298), .A2(crash_dump_o_65_), .ZN(n2297) );
NAND2_X1 U25991 ( .A1(n11459), .A2(n19960), .ZN(n2298) );
NAND2_X1 U25992 ( .A1(n5714), .A2(n10280), .ZN(n5671) );
NAND2_X1 U25993 ( .A1(n11320), .A2(n10281), .ZN(n10280) );
NAND2_X1 U25994 ( .A1(n11329), .A2(n15858), .ZN(n10281) );
NAND2_X1 U25995 ( .A1(n11290), .A2(n11289), .ZN(n4927) );
NAND2_X1 U25996 ( .A1(n10147), .A2(n10146), .ZN(n10133) );
NOR2_X1 U25997 ( .A1(n10151), .A2(n1687), .ZN(n10147) );
NOR2_X1 U25998 ( .A1(n11327), .A2(n10144), .ZN(n10151) );
OR2_X1 U25999 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_1), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_0), .ZN(n22103) );
OR2_X1 U26000 ( .A1(n22103), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_2), .ZN(n22105) );
OR2_X1 U26001 ( .A1(n22105), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_3), .ZN(n22107) );
NAND2_X1 U26002 ( .A1(n11519), .A2(id_stage_i_controller_i_do_single_step_q), .ZN(n5131) );
AND2_X1 U26003 ( .A1(n10081), .A2(n10082), .ZN(n15773) );
NOR2_X1 U26004 ( .A1(n10266), .A2(n10267), .ZN(n10081) );
NOR2_X1 U26005 ( .A1(n1440), .A2(n10083), .ZN(n10082) );
NAND2_X1 U26006 ( .A1(n20912), .A2(n11502), .ZN(n10267) );
NOR2_X1 U26007 ( .A1(n11472), .A2(n3019), .ZN(n15752) );
NAND2_X1 U26008 ( .A1(n2192), .A2(crash_dump_o_65_), .ZN(n2191) );
NAND2_X1 U26009 ( .A1(n2193), .A2(n2194), .ZN(n2192) );
NAND2_X1 U26010 ( .A1(n11459), .A2(instr_rdata_i_6_), .ZN(n2194) );
NAND2_X1 U26011 ( .A1(n15803), .A2(n16045), .ZN(n2193) );
NAND2_X1 U26012 ( .A1(n2254), .A2(crash_dump_o_65_), .ZN(n2253) );
NAND2_X1 U26013 ( .A1(n2255), .A2(n2256), .ZN(n2254) );
NAND2_X1 U26014 ( .A1(n11459), .A2(instr_rdata_i_3_), .ZN(n2256) );
NAND2_X1 U26015 ( .A1(n15803), .A2(n16046), .ZN(n2255) );
AND2_X1 U26016 ( .A1(n15925), .A2(n1583), .ZN(n1527) );
NAND2_X1 U26017 ( .A1(n11298), .A2(n11296), .ZN(n1583) );
NOR2_X1 U26018 ( .A1(n6756), .A2(n6757), .ZN(n6754) );
NOR2_X1 U26019 ( .A1(n11354), .A2(n6712), .ZN(n6756) );
NOR2_X1 U26020 ( .A1(n19801), .A2(n6711), .ZN(n6757) );
NOR2_X1 U26021 ( .A1(n6778), .A2(n6779), .ZN(n6776) );
NOR2_X1 U26022 ( .A1(n11350), .A2(n6712), .ZN(n6778) );
NOR2_X1 U26023 ( .A1(n19805), .A2(n6711), .ZN(n6779) );
NOR2_X1 U26024 ( .A1(n6810), .A2(n6811), .ZN(n6808) );
NOR2_X1 U26025 ( .A1(n11348), .A2(n6712), .ZN(n6810) );
NOR2_X1 U26026 ( .A1(n19807), .A2(n6711), .ZN(n6811) );
NOR2_X1 U26027 ( .A1(n6912), .A2(n6913), .ZN(n6910) );
NOR2_X1 U26028 ( .A1(n11346), .A2(n6712), .ZN(n6912) );
NOR2_X1 U26029 ( .A1(n19809), .A2(n6711), .ZN(n6913) );
NOR2_X1 U26030 ( .A1(n6989), .A2(n6990), .ZN(n6987) );
NOR2_X1 U26031 ( .A1(n11366), .A2(n6712), .ZN(n6989) );
NOR2_X1 U26032 ( .A1(n19787), .A2(n6711), .ZN(n6990) );
NOR2_X1 U26033 ( .A1(n6999), .A2(n7000), .ZN(n6997) );
NOR2_X1 U26034 ( .A1(n11364), .A2(n6712), .ZN(n6999) );
NOR2_X1 U26035 ( .A1(n19789), .A2(n6711), .ZN(n7000) );
NOR2_X1 U26036 ( .A1(n7020), .A2(n7021), .ZN(n7017) );
NOR2_X1 U26037 ( .A1(n11374), .A2(n6712), .ZN(n7020) );
NOR2_X1 U26038 ( .A1(n19811), .A2(n6711), .ZN(n7021) );
NOR2_X1 U26039 ( .A1(n6959), .A2(n6960), .ZN(n6957) );
NOR2_X1 U26040 ( .A1(n11372), .A2(n6712), .ZN(n6959) );
NOR2_X1 U26041 ( .A1(n19781), .A2(n6711), .ZN(n6960) );
NOR2_X1 U26042 ( .A1(n6969), .A2(n6970), .ZN(n6967) );
NOR2_X1 U26043 ( .A1(n11370), .A2(n6712), .ZN(n6969) );
NOR2_X1 U26044 ( .A1(n19783), .A2(n6711), .ZN(n6970) );
NOR2_X1 U26045 ( .A1(n6979), .A2(n6980), .ZN(n6977) );
NOR2_X1 U26046 ( .A1(n11368), .A2(n6712), .ZN(n6979) );
NOR2_X1 U26047 ( .A1(n19785), .A2(n6711), .ZN(n6980) );
NOR2_X1 U26048 ( .A1(n7009), .A2(n7010), .ZN(n7007) );
NOR2_X1 U26049 ( .A1(n11463), .A2(n6712), .ZN(n7009) );
NOR2_X1 U26050 ( .A1(n19791), .A2(n6711), .ZN(n7010) );
NOR2_X1 U26051 ( .A1(n6709), .A2(n6710), .ZN(n6706) );
NOR2_X1 U26052 ( .A1(n11362), .A2(n6712), .ZN(n6709) );
NOR2_X1 U26053 ( .A1(n19793), .A2(n6711), .ZN(n6710) );
NOR2_X1 U26054 ( .A1(n6724), .A2(n6725), .ZN(n6722) );
NOR2_X1 U26055 ( .A1(n11360), .A2(n6712), .ZN(n6724) );
NOR2_X1 U26056 ( .A1(n19795), .A2(n6711), .ZN(n6725) );
NOR2_X1 U26057 ( .A1(n6745), .A2(n6746), .ZN(n6743) );
NOR2_X1 U26058 ( .A1(n11356), .A2(n6712), .ZN(n6745) );
NOR2_X1 U26059 ( .A1(n19799), .A2(n6711), .ZN(n6746) );
NOR2_X1 U26060 ( .A1(n6767), .A2(n6768), .ZN(n6765) );
NOR2_X1 U26061 ( .A1(n11352), .A2(n6712), .ZN(n6767) );
NOR2_X1 U26062 ( .A1(n19803), .A2(n6711), .ZN(n6768) );
NOR2_X1 U26063 ( .A1(n6734), .A2(n6735), .ZN(n6732) );
NOR2_X1 U26064 ( .A1(n11358), .A2(n6712), .ZN(n6734) );
NOR2_X1 U26065 ( .A1(n19797), .A2(n6711), .ZN(n6735) );
AND2_X1 U26066 ( .A1(n10071), .A2(n10072), .ZN(n10066) );
NOR2_X1 U26067 ( .A1(n11320), .A2(n10074), .ZN(n10071) );
NOR2_X1 U26068 ( .A1(rf_raddr_a_o_2_), .A2(n10073), .ZN(n10072) );
NAND2_X1 U26069 ( .A1(n15890), .A2(n15809), .ZN(n10074) );
NAND2_X1 U26070 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N219), .A2(n5065), .ZN(n5064) );
NAND2_X1 U26071 ( .A1(n11285), .A2(n21006), .ZN(n5065) );
NAND2_X1 U26072 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N219), .A2(n5045), .ZN(n5044) );
NAND2_X1 U26073 ( .A1(n11262), .A2(n21006), .ZN(n5045) );
INV_X1 U26074 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_31_), .ZN(n20080) );
NAND2_X1 U26075 ( .A1(n11090), .A2(n1500), .ZN(n1452) );
NAND2_X1 U26076 ( .A1(n1501), .A2(n1502), .ZN(n1500) );
NAND2_X1 U26077 ( .A1(n20997), .A2(data_rvalid_i), .ZN(n1502) );
NAND2_X1 U26078 ( .A1(n10065), .A2(n20937), .ZN(n8557) );
NOR2_X1 U26079 ( .A1(n11320), .A2(n10066), .ZN(n10065) );
AND2_X1 U26080 ( .A1(n10426), .A2(n10427), .ZN(n5251) );
NOR2_X1 U26081 ( .A1(rf_raddr_b_o_1_), .A2(n10431), .ZN(n10426) );
NOR2_X1 U26082 ( .A1(n11338), .A2(n10428), .ZN(n10427) );
NAND2_X1 U26083 ( .A1(n20969), .A2(n10287), .ZN(n10431) );
NOR2_X1 U26084 ( .A1(n3019), .A2(n3705), .ZN(n15748) );
NOR2_X1 U26085 ( .A1(n16132), .A2(n3707), .ZN(n3705) );
NAND2_X1 U26086 ( .A1(n3708), .A2(n3709), .ZN(n3707) );
NAND2_X1 U26087 ( .A1(n19873), .A2(n11458), .ZN(n3129) );
NAND2_X1 U26088 ( .A1(n19874), .A2(n11459), .ZN(n3262) );
NOR2_X1 U26089 ( .A1(n11485), .A2(n2532), .ZN(n2530) );
NOR2_X1 U26090 ( .A1(instr_rdata_i_14_), .A2(n15803), .ZN(n2532) );
NAND2_X1 U26091 ( .A1(n11023), .A2(n19971), .ZN(n15273) );
AND2_X1 U26092 ( .A1(n10472), .A2(n11515), .ZN(n10464) );
NOR2_X1 U26093 ( .A1(n11514), .A2(n11516), .ZN(n10472) );
NOR2_X1 U26094 ( .A1(n21486), .A2(n21485), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_3) );
NOR2_X1 U26095 ( .A1(crash_dump_o_67_), .A2(n21491), .ZN(n21485) );
NOR2_X1 U26096 ( .A1(n11030), .A2(n6561), .ZN(n15280) );
NOR2_X1 U26097 ( .A1(n11029), .A2(n6561), .ZN(n15279) );
NOR2_X1 U26098 ( .A1(n11028), .A2(n6561), .ZN(n15278) );
NOR2_X1 U26099 ( .A1(n11027), .A2(n6561), .ZN(n15277) );
NOR2_X1 U26100 ( .A1(n11026), .A2(n6561), .ZN(n15276) );
NOR2_X1 U26101 ( .A1(n11025), .A2(n6561), .ZN(n15275) );
NOR2_X1 U26102 ( .A1(n11024), .A2(n6561), .ZN(n15274) );
AND2_X1 U26103 ( .A1(n11517), .A2(n8074), .ZN(n8070) );
NAND2_X1 U26104 ( .A1(n10765), .A2(n10351), .ZN(n5271) );
OR2_X1 U26105 ( .A1(n10266), .A2(n10276), .ZN(n10351) );
NAND2_X1 U26106 ( .A1(n10456), .A2(n10457), .ZN(n5269) );
NOR2_X1 U26107 ( .A1(n11340), .A2(rf_raddr_b_o_2_), .ZN(n10456) );
NOR2_X1 U26108 ( .A1(n11336), .A2(n10458), .ZN(n10457) );
OR2_X1 U26109 ( .A1(n11325), .A2(n11311), .ZN(n10458) );
AND2_X1 U26110 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_4), .A2(n11253), .ZN(n22087) );
AND2_X1 U26111 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_3), .ZN(n22091) );
NAND2_X1 U26112 ( .A1(n5713), .A2(n5714), .ZN(n5532) );
NOR2_X1 U26113 ( .A1(n11320), .A2(n15858), .ZN(n5713) );
NAND2_X1 U26114 ( .A1(n20931), .A2(n10349), .ZN(n10321) );
NAND2_X1 U26115 ( .A1(n10350), .A2(n10766), .ZN(n10349) );
AND2_X1 U26116 ( .A1(n5271), .A2(n20984), .ZN(n10350) );
NAND2_X1 U26117 ( .A1(n2573), .A2(n2574), .ZN(n2570) );
NOR2_X1 U26118 ( .A1(n2578), .A2(n2579), .ZN(n2573) );
NOR2_X1 U26119 ( .A1(n2575), .A2(n2576), .ZN(n2574) );
NOR2_X1 U26120 ( .A1(n11386), .A2(n16448), .ZN(n2579) );
NAND2_X1 U26121 ( .A1(n2602), .A2(n2603), .ZN(n2599) );
NOR2_X1 U26122 ( .A1(n2607), .A2(n2608), .ZN(n2602) );
NOR2_X1 U26123 ( .A1(n2604), .A2(n2605), .ZN(n2603) );
NOR2_X1 U26124 ( .A1(n11385), .A2(n2169), .ZN(n2608) );
NAND2_X1 U26125 ( .A1(crash_dump_o_126_), .A2(n20898), .ZN(n21595) );
INV_X1 U26126 ( .A(n21594), .ZN(n20898) );
NAND2_X1 U26127 ( .A1(n7713), .A2(n7712), .ZN(n7662) );
NOR2_X1 U26128 ( .A1(n10546), .A2(n20923), .ZN(n7713) );
NOR2_X1 U26129 ( .A1(n11464), .A2(n16450), .ZN(n15743) );
INV_X1 U26130 ( .A(instr_rdata_i_17_), .ZN(n19944) );
NAND2_X1 U26131 ( .A1(n11313), .A2(n10374), .ZN(n10446) );
NAND2_X1 U26132 ( .A1(n7003), .A2(n7004), .ZN(n7002) );
NAND2_X1 U26133 ( .A1(n20875), .A2(rf_waddr_wb_o_4_), .ZN(n7003) );
NAND2_X1 U26134 ( .A1(n20876), .A2(crash_dump_o_43_), .ZN(n7004) );
NAND2_X1 U26135 ( .A1(n6963), .A2(n6964), .ZN(n6962) );
NAND2_X1 U26136 ( .A1(n20875), .A2(rf_raddr_a_o_0_), .ZN(n6963) );
NAND2_X1 U26137 ( .A1(n20876), .A2(crash_dump_o_47_), .ZN(n6964) );
NAND2_X1 U26138 ( .A1(n7013), .A2(n7014), .ZN(n7012) );
NAND2_X1 U26139 ( .A1(n20875), .A2(rf_waddr_wb_o_3_), .ZN(n7013) );
NAND2_X1 U26140 ( .A1(n20876), .A2(crash_dump_o_42_), .ZN(n7014) );
NAND2_X1 U26141 ( .A1(n6715), .A2(n6716), .ZN(n6714) );
NAND2_X1 U26142 ( .A1(n20875), .A2(rf_waddr_wb_o_2_), .ZN(n6715) );
NAND2_X1 U26143 ( .A1(n20876), .A2(crash_dump_o_41_), .ZN(n6716) );
NAND2_X1 U26144 ( .A1(n6728), .A2(n6729), .ZN(n6727) );
NAND2_X1 U26145 ( .A1(n20875), .A2(rf_waddr_wb_o_1_), .ZN(n6728) );
NAND2_X1 U26146 ( .A1(n20876), .A2(crash_dump_o_40_), .ZN(n6729) );
NAND2_X1 U26147 ( .A1(n6739), .A2(n6740), .ZN(n6738) );
NAND2_X1 U26148 ( .A1(n20875), .A2(rf_waddr_wb_o_0_), .ZN(n6739) );
NAND2_X1 U26149 ( .A1(n20876), .A2(crash_dump_o_39_), .ZN(n6740) );
NAND2_X1 U26150 ( .A1(n4753), .A2(n4754), .ZN(n4752) );
NAND2_X1 U26151 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_2), .ZN(n4753) );
NAND2_X1 U26152 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_18), .A2(n4275), .ZN(n4754) );
NAND2_X1 U26153 ( .A1(n4693), .A2(n4694), .ZN(n4692) );
NAND2_X1 U26154 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_4), .ZN(n4693) );
NAND2_X1 U26155 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_20), .A2(n4275), .ZN(n4694) );
NAND2_X1 U26156 ( .A1(n4672), .A2(n4673), .ZN(n4671) );
NAND2_X1 U26157 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_5), .ZN(n4672) );
NAND2_X1 U26158 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_21), .A2(n4275), .ZN(n4673) );
NAND2_X1 U26159 ( .A1(n4630), .A2(n4631), .ZN(n4629) );
NAND2_X1 U26160 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_7), .ZN(n4630) );
NAND2_X1 U26161 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_23), .A2(n4275), .ZN(n4631) );
NAND2_X1 U26162 ( .A1(n4440), .A2(n4441), .ZN(n4439) );
NAND2_X1 U26163 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_15), .ZN(n4440) );
NAND2_X1 U26164 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_31), .A2(n4275), .ZN(n4441) );
NAND2_X1 U26165 ( .A1(n4795), .A2(n4796), .ZN(n4794) );
NAND2_X1 U26166 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_0), .ZN(n4795) );
NAND2_X1 U26167 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_16), .A2(n4275), .ZN(n4796) );
NAND2_X1 U26168 ( .A1(n4774), .A2(n4775), .ZN(n4773) );
NAND2_X1 U26169 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_1), .ZN(n4774) );
NAND2_X1 U26170 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_17), .A2(n16423), .ZN(n4775) );
NAND2_X1 U26171 ( .A1(n4732), .A2(n4733), .ZN(n4731) );
NAND2_X1 U26172 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_3), .ZN(n4732) );
NAND2_X1 U26173 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_19), .A2(n16423), .ZN(n4733) );
NAND2_X1 U26174 ( .A1(n4651), .A2(n4652), .ZN(n4650) );
NAND2_X1 U26175 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_6), .ZN(n4651) );
NAND2_X1 U26176 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_22), .A2(n16423), .ZN(n4652) );
NAND2_X1 U26177 ( .A1(n4609), .A2(n4610), .ZN(n4608) );
NAND2_X1 U26178 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_8), .ZN(n4609) );
NAND2_X1 U26179 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_24), .A2(n16423), .ZN(n4610) );
NAND2_X1 U26180 ( .A1(n4588), .A2(n4589), .ZN(n4587) );
NAND2_X1 U26181 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_9), .ZN(n4588) );
NAND2_X1 U26182 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_25), .A2(n16423), .ZN(n4589) );
NAND2_X1 U26183 ( .A1(n4567), .A2(n4568), .ZN(n4566) );
NAND2_X1 U26184 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_10), .ZN(n4567) );
NAND2_X1 U26185 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_26), .A2(n4275), .ZN(n4568) );
NAND2_X1 U26186 ( .A1(n4546), .A2(n4547), .ZN(n4545) );
NAND2_X1 U26187 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_11), .ZN(n4546) );
NAND2_X1 U26188 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_27), .A2(n16423), .ZN(n4547) );
NAND2_X1 U26189 ( .A1(n4525), .A2(n4526), .ZN(n4524) );
NAND2_X1 U26190 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_12), .ZN(n4525) );
NAND2_X1 U26191 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_28), .A2(n16423), .ZN(n4526) );
NAND2_X1 U26192 ( .A1(n4504), .A2(n4505), .ZN(n4503) );
NAND2_X1 U26193 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_13), .ZN(n4504) );
NAND2_X1 U26194 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_29), .A2(n16423), .ZN(n4505) );
NAND2_X1 U26195 ( .A1(n4464), .A2(n4465), .ZN(n4463) );
NAND2_X1 U26196 ( .A1(n20907), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_14), .ZN(n4464) );
NAND2_X1 U26197 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_30), .A2(n4275), .ZN(n4465) );
NAND2_X1 U26198 ( .A1(data_gnt_i), .A2(n1576), .ZN(n1601) );
NAND2_X1 U26199 ( .A1(n2751), .A2(n2752), .ZN(n2750) );
NAND2_X1 U26200 ( .A1(n11423), .A2(n15803), .ZN(n2751) );
NAND2_X1 U26201 ( .A1(n2753), .A2(n11459), .ZN(n2752) );
NAND2_X1 U26202 ( .A1(n10363), .A2(n15876), .ZN(n10361) );
NAND2_X1 U26203 ( .A1(n10364), .A2(n10365), .ZN(n10363) );
NAND2_X1 U26204 ( .A1(n10368), .A2(n11320), .ZN(n10364) );
NAND2_X1 U26205 ( .A1(n10366), .A2(n10367), .ZN(n10365) );
NAND2_X1 U26206 ( .A1(n8885), .A2(n8886), .ZN(n8452) );
NAND2_X1 U26207 ( .A1(n8310), .A2(n20852), .ZN(n8886) );
NAND2_X1 U26208 ( .A1(n11509), .A2(n8883), .ZN(n8885) );
NAND2_X1 U26209 ( .A1(n5019), .A2(n21010), .ZN(n5018) );
NAND2_X1 U26210 ( .A1(n11274), .A2(n5010), .ZN(n5019) );
NAND2_X1 U26211 ( .A1(n5077), .A2(n5078), .ZN(n5072) );
NAND2_X1 U26212 ( .A1(n11257), .A2(n5011), .ZN(n5078) );
NOR2_X1 U26213 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N219), .A2(n5079), .ZN(n5077) );
NOR2_X1 U26214 ( .A1(n21007), .A2(n16120), .ZN(n5079) );
NAND2_X1 U26215 ( .A1(n5056), .A2(n5057), .ZN(n5052) );
NAND2_X1 U26216 ( .A1(n11287), .A2(n5011), .ZN(n5057) );
NOR2_X1 U26217 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N219), .A2(n5058), .ZN(n5056) );
NOR2_X1 U26218 ( .A1(n21007), .A2(n16121), .ZN(n5058) );
NAND2_X1 U26219 ( .A1(n5008), .A2(n5009), .ZN(n5002) );
NAND2_X1 U26220 ( .A1(n11265), .A2(n5010), .ZN(n5009) );
NAND2_X1 U26221 ( .A1(n11264), .A2(n5011), .ZN(n5008) );
NAND2_X1 U26222 ( .A1(n10209), .A2(n10201), .ZN(n10208) );
NAND2_X1 U26223 ( .A1(n20981), .A2(n10211), .ZN(n10209) );
NAND2_X1 U26224 ( .A1(n10212), .A2(n10213), .ZN(n10211) );
NAND2_X1 U26225 ( .A1(n20946), .A2(n11328), .ZN(n10212) );
NAND2_X1 U26226 ( .A1(crash_dump_o_117_), .A2(n21563), .ZN(n21558) );
NAND2_X1 U26227 ( .A1(crash_dump_o_123_), .A2(n21584), .ZN(n21579) );
NAND2_X1 U26228 ( .A1(crash_dump_o_121_), .A2(n21577), .ZN(n21572) );
NAND2_X1 U26229 ( .A1(crash_dump_o_119_), .A2(n21570), .ZN(n21565) );
NAND2_X1 U26230 ( .A1(crash_dump_o_115_), .A2(n21556), .ZN(n21549) );
NAND2_X1 U26231 ( .A1(crash_dump_o_113_), .A2(n21547), .ZN(n21542) );
NAND2_X1 U26232 ( .A1(n2551), .A2(n2552), .ZN(n2550) );
NAND2_X1 U26233 ( .A1(n11404), .A2(n15803), .ZN(n2552) );
NOR2_X1 U26234 ( .A1(n11485), .A2(n2553), .ZN(n2551) );
NOR2_X1 U26235 ( .A1(instr_rdata_i_13_), .A2(n15803), .ZN(n2553) );
NAND2_X1 U26236 ( .A1(n5030), .A2(n5031), .ZN(n5029) );
NAND2_X1 U26237 ( .A1(n11278), .A2(n5010), .ZN(n5031) );
NAND2_X1 U26238 ( .A1(n11277), .A2(n5011), .ZN(n5030) );
NAND2_X1 U26239 ( .A1(n11484), .A2(n20938), .ZN(n10398) );
NAND2_X1 U26240 ( .A1(n11263), .A2(n21008), .ZN(n5047) );
NAND2_X1 U26241 ( .A1(n11267), .A2(n21008), .ZN(n5005) );
NAND2_X1 U26242 ( .A1(n10375), .A2(n10376), .ZN(n10355) );
OR2_X1 U26243 ( .A1(n1442), .A2(n10377), .ZN(n10376) );
NOR2_X1 U26244 ( .A1(n10378), .A2(n10379), .ZN(n10375) );
NOR2_X1 U26245 ( .A1(n11504), .A2(n10380), .ZN(n10379) );
NAND2_X1 U26246 ( .A1(crash_dump_o_125_), .A2(n21591), .ZN(n21586) );
NAND2_X1 U26247 ( .A1(n5066), .A2(n5067), .ZN(n5063) );
NAND2_X1 U26248 ( .A1(n11286), .A2(n21008), .ZN(n5067) );
NOR2_X1 U26249 ( .A1(n5068), .A2(n5069), .ZN(n5066) );
NOR2_X1 U26250 ( .A1(n21009), .A2(n16122), .ZN(n5069) );
NAND2_X1 U26251 ( .A1(n11266), .A2(n21006), .ZN(n5004) );
NAND2_X1 U26252 ( .A1(n10240), .A2(n10241), .ZN(n10239) );
NAND2_X1 U26253 ( .A1(n10245), .A2(n11322), .ZN(n10240) );
NAND2_X1 U26254 ( .A1(n10242), .A2(n20978), .ZN(n10241) );
NOR2_X1 U26255 ( .A1(n11317), .A2(n11327), .ZN(n10245) );
NAND2_X1 U26256 ( .A1(n5074), .A2(n5075), .ZN(n5073) );
NAND2_X1 U26257 ( .A1(n11279), .A2(n21006), .ZN(n5074) );
NAND2_X1 U26258 ( .A1(n11282), .A2(n21008), .ZN(n5075) );
NAND2_X1 U26259 ( .A1(n5054), .A2(n5055), .ZN(n5053) );
NAND2_X1 U26260 ( .A1(n11258), .A2(n21006), .ZN(n5054) );
NAND2_X1 U26261 ( .A1(n11259), .A2(n21008), .ZN(n5055) );
NAND2_X1 U26262 ( .A1(crash_dump_o_126_), .A2(n21594), .ZN(n21592) );
INV_X1 U26263 ( .A(n25267), .ZN(n20028) );
NAND2_X1 U26264 ( .A1(instr_rdata_i_30_), .A2(n16447), .ZN(n2528) );
NAND2_X1 U26265 ( .A1(instr_rdata_i_21_), .A2(n16447), .ZN(n2212) );
NAND2_X1 U26266 ( .A1(instr_rdata_i_24_), .A2(n16447), .ZN(n2121) );
NAND2_X1 U26267 ( .A1(n10401), .A2(n15884), .ZN(n10400) );
NAND2_X1 U26268 ( .A1(n20977), .A2(n10403), .ZN(n10401) );
INV_X1 U26269 ( .A(n1442), .ZN(n20977) );
NAND2_X1 U26270 ( .A1(n11504), .A2(n15804), .ZN(n10403) );
NAND2_X1 U26271 ( .A1(crash_dump_o_122_), .A2(n21574), .ZN(n21575) );
NAND2_X1 U26272 ( .A1(crash_dump_o_120_), .A2(n21567), .ZN(n21568) );
NAND2_X1 U26273 ( .A1(crash_dump_o_118_), .A2(n21560), .ZN(n21561) );
NAND2_X1 U26274 ( .A1(crash_dump_o_116_), .A2(n21553), .ZN(n21554) );
NAND2_X1 U26275 ( .A1(crash_dump_o_114_), .A2(n21544), .ZN(n21545) );
NAND2_X1 U26276 ( .A1(crash_dump_o_112_), .A2(n21537), .ZN(n21538) );
NAND2_X1 U26277 ( .A1(crash_dump_o_124_), .A2(n21581), .ZN(n21582) );
NAND2_X1 U26278 ( .A1(n10084), .A2(n15917), .ZN(n10083) );
NAND2_X1 U26279 ( .A1(n11292), .A2(n1412), .ZN(n10084) );
NAND2_X1 U26280 ( .A1(n10440), .A2(n10441), .ZN(n10416) );
NOR2_X1 U26281 ( .A1(rf_raddr_a_o_4_), .A2(n10444), .ZN(n10440) );
NOR2_X1 U26282 ( .A1(rf_waddr_wb_o_2_), .A2(n10442), .ZN(n10441) );
NAND2_X1 U26283 ( .A1(n16123), .A2(n15828), .ZN(n10444) );
NAND2_X1 U26284 ( .A1(instr_rdata_i_22_), .A2(n16447), .ZN(n2190) );
NAND2_X1 U26285 ( .A1(instr_rdata_i_19_), .A2(n16447), .ZN(n2252) );
NAND2_X1 U26286 ( .A1(n11475), .A2(n11515), .ZN(n10462) );
NAND2_X1 U26287 ( .A1(n10418), .A2(n10419), .ZN(n10417) );
NOR2_X1 U26288 ( .A1(n5258), .A2(n10421), .ZN(n10418) );
NOR2_X1 U26289 ( .A1(rf_raddr_a_o_1_), .A2(n10420), .ZN(n10419) );
NAND2_X1 U26290 ( .A1(n10422), .A2(n15890), .ZN(n10421) );
NAND2_X1 U26291 ( .A1(n5263), .A2(n5264), .ZN(n5262) );
NOR2_X1 U26292 ( .A1(rf_raddr_b_o_0_), .A2(n5266), .ZN(n5264) );
NAND2_X1 U26293 ( .A1(n11336), .A2(n5267), .ZN(n5266) );
NAND2_X1 U26294 ( .A1(n11503), .A2(n11501), .ZN(n10362) );
NAND2_X1 U26295 ( .A1(instr_rdata_i_0_), .A2(n11460), .ZN(n3606) );
NAND2_X1 U26296 ( .A1(n11255), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_0), .ZN(n5562) );
NAND2_X1 U26297 ( .A1(crash_dump_o_127_), .A2(n21595), .ZN(n21596) );
NAND2_X1 U26298 ( .A1(n2746), .A2(n11485), .ZN(n2745) );
OR2_X1 U26299 ( .A1(n1446), .A2(instr_gnt_i), .ZN(n2897) );
NAND2_X1 U26300 ( .A1(n11290), .A2(n4965), .ZN(n4964) );
NAND2_X1 U26301 ( .A1(n4966), .A2(n4967), .ZN(n4965) );
NAND2_X1 U26302 ( .A1(n21000), .A2(rf_rdata_a_ecc_i_0_), .ZN(n4966) );
NAND2_X1 U26303 ( .A1(n4968), .A2(n20919), .ZN(n4967) );
AND2_X1 U26304 ( .A1(n5239), .A2(n4056), .ZN(n15564) );
NAND2_X1 U26305 ( .A1(n5240), .A2(n5241), .ZN(n5239) );
OR2_X1 U26306 ( .A1(n5242), .A2(n11519), .ZN(n5241) );
NOR2_X1 U26307 ( .A1(n5243), .A2(n5244), .ZN(n5240) );
NAND2_X1 U26308 ( .A1(n11459), .A2(n19946), .ZN(n2505) );
NAND2_X1 U26309 ( .A1(n21605), .A2(n21604), .ZN(id_stage_i_controller_i_N262) );
OR2_X1 U26310 ( .A1(n21606), .A2(crash_dump_o_101_), .ZN(n21605) );
NAND2_X1 U26311 ( .A1(crash_dump_o_101_), .A2(n21606), .ZN(n21604) );
NAND2_X1 U26312 ( .A1(n21599), .A2(n21598), .ZN(id_stage_i_controller_i_N260) );
OR2_X1 U26313 ( .A1(n21600), .A2(crash_dump_o_99_), .ZN(n21599) );
NAND2_X1 U26314 ( .A1(crash_dump_o_99_), .A2(n21600), .ZN(n21598) );
NAND2_X1 U26315 ( .A1(n21522), .A2(n21521), .ZN(id_stage_i_controller_i_N268) );
OR2_X1 U26316 ( .A1(n21526), .A2(crash_dump_o_107_), .ZN(n21522) );
NAND2_X1 U26317 ( .A1(crash_dump_o_107_), .A2(n21526), .ZN(n21521) );
NAND2_X1 U26318 ( .A1(n21536), .A2(n21535), .ZN(id_stage_i_controller_i_N272) );
OR2_X1 U26319 ( .A1(n21540), .A2(crash_dump_o_111_), .ZN(n21536) );
NAND2_X1 U26320 ( .A1(crash_dump_o_111_), .A2(n21540), .ZN(n21535) );
NAND2_X1 U26321 ( .A1(n21529), .A2(n21528), .ZN(id_stage_i_controller_i_N270) );
OR2_X1 U26322 ( .A1(n21533), .A2(crash_dump_o_109_), .ZN(n21529) );
NAND2_X1 U26323 ( .A1(crash_dump_o_109_), .A2(n21533), .ZN(n21528) );
NAND2_X1 U26324 ( .A1(n21611), .A2(n21610), .ZN(id_stage_i_controller_i_N264) );
OR2_X1 U26325 ( .A1(n21612), .A2(crash_dump_o_103_), .ZN(n21611) );
NAND2_X1 U26326 ( .A1(crash_dump_o_103_), .A2(n21612), .ZN(n21610) );
NAND2_X1 U26327 ( .A1(n21618), .A2(n21617), .ZN(id_stage_i_controller_i_N266) );
OR2_X1 U26328 ( .A1(n21616), .A2(crash_dump_o_105_), .ZN(n21618) );
NAND2_X1 U26329 ( .A1(crash_dump_o_105_), .A2(n21616), .ZN(n21617) );
NAND2_X1 U26330 ( .A1(n10393), .A2(n10394), .ZN(n10392) );
NOR2_X1 U26331 ( .A1(n15807), .A2(n15879), .ZN(n10393) );
NOR2_X1 U26332 ( .A1(n10395), .A2(n10396), .ZN(n10394) );
NOR2_X1 U26333 ( .A1(n11313), .A2(n15805), .ZN(n10396) );
NAND2_X1 U26334 ( .A1(n21552), .A2(n21551), .ZN(id_stage_i_controller_i_N258) );
NAND2_X1 U26335 ( .A1(crash_dump_o_97_), .A2(n15928), .ZN(n21552) );
NAND2_X1 U26336 ( .A1(instr_fetch_err_plus2), .A2(n11465), .ZN(n21551) );
INV_X1 U26337 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N67), .ZN(n20024) );
NAND2_X1 U26338 ( .A1(n20954), .A2(rf_waddr_wb_o_0_), .ZN(n10511) );
NAND2_X1 U26339 ( .A1(n5082), .A2(n11289), .ZN(n5081) );
NOR2_X1 U26340 ( .A1(n11281), .A2(n11290), .ZN(n5082) );
NAND2_X1 U26341 ( .A1(n20902), .A2(instr_rdata_i_5_), .ZN(n2215) );
NAND2_X1 U26342 ( .A1(n20902), .A2(instr_rdata_i_8_), .ZN(n2126) );
NAND2_X1 U26343 ( .A1(n21525), .A2(n21524), .ZN(id_stage_i_controller_i_N269) );
OR2_X1 U26344 ( .A1(n21523), .A2(crash_dump_o_108_), .ZN(n21525) );
NAND2_X1 U26345 ( .A1(crash_dump_o_108_), .A2(n21523), .ZN(n21524) );
OR2_X1 U26346 ( .A1(n11307), .A2(n21526), .ZN(n21523) );
NAND2_X1 U26347 ( .A1(n21532), .A2(n21531), .ZN(id_stage_i_controller_i_N271) );
OR2_X1 U26348 ( .A1(n21530), .A2(crash_dump_o_110_), .ZN(n21532) );
NAND2_X1 U26349 ( .A1(crash_dump_o_110_), .A2(n21530), .ZN(n21531) );
OR2_X1 U26350 ( .A1(n10788), .A2(n21533), .ZN(n21530) );
NAND2_X1 U26351 ( .A1(n21615), .A2(n21614), .ZN(id_stage_i_controller_i_N265) );
OR2_X1 U26352 ( .A1(n21613), .A2(crash_dump_o_104_), .ZN(n21615) );
NAND2_X1 U26353 ( .A1(crash_dump_o_104_), .A2(n21613), .ZN(n21614) );
OR2_X1 U26354 ( .A1(n10680), .A2(n21612), .ZN(n21613) );
NAND2_X1 U26355 ( .A1(n21609), .A2(n21608), .ZN(id_stage_i_controller_i_N263) );
OR2_X1 U26356 ( .A1(n21607), .A2(crash_dump_o_102_), .ZN(n21609) );
NAND2_X1 U26357 ( .A1(crash_dump_o_102_), .A2(n21607), .ZN(n21608) );
OR2_X1 U26358 ( .A1(n11466), .A2(n21606), .ZN(n21607) );
NAND2_X1 U26359 ( .A1(n21603), .A2(n21602), .ZN(id_stage_i_controller_i_N261) );
OR2_X1 U26360 ( .A1(n21601), .A2(crash_dump_o_100_), .ZN(n21603) );
NAND2_X1 U26361 ( .A1(crash_dump_o_100_), .A2(n21601), .ZN(n21602) );
OR2_X1 U26362 ( .A1(n10670), .A2(n21600), .ZN(n21601) );
NAND2_X1 U26363 ( .A1(n21519), .A2(n21518), .ZN(id_stage_i_controller_i_N267) );
OR2_X1 U26364 ( .A1(n21517), .A2(crash_dump_o_106_), .ZN(n21519) );
NAND2_X1 U26365 ( .A1(crash_dump_o_106_), .A2(n21517), .ZN(n21518) );
OR2_X1 U26366 ( .A1(n21616), .A2(n10745), .ZN(n21517) );
AND2_X1 U26367 ( .A1(n3050), .A2(n11460), .ZN(n3582) );
AND2_X1 U26368 ( .A1(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_1), .A2(n16432), .ZN(n3495) );
NOR2_X1 U26369 ( .A1(n21405), .A2(n21446), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_1) );
NOR2_X1 U26370 ( .A1(crash_dump_o_65_), .A2(n19938), .ZN(n21405) );
AND2_X1 U26371 ( .A1(n10516), .A2(n11328), .ZN(n10529) );
AND2_X1 U26372 ( .A1(n10102), .A2(n11328), .ZN(n10101) );
INV_X1 U26373 ( .A(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N68), .ZN(n20025) );
OR2_X1 U26374 ( .A1(n20931), .A2(n11306), .ZN(n3971) );
OR2_X1 U26375 ( .A1(n20931), .A2(n10840), .ZN(n3915) );
OR2_X1 U26376 ( .A1(n20931), .A2(n10887), .ZN(n3870) );
OR2_X1 U26377 ( .A1(n20931), .A2(n10947), .ZN(n3814) );
OR2_X1 U26378 ( .A1(n20931), .A2(n10977), .ZN(n3791) );
OR2_X1 U26379 ( .A1(n20931), .A2(n10634), .ZN(n3779) );
OR2_X1 U26380 ( .A1(n21563), .A2(crash_dump_o_117_), .ZN(n21559) );
OR2_X1 U26381 ( .A1(n21584), .A2(crash_dump_o_123_), .ZN(n21580) );
OR2_X1 U26382 ( .A1(n21577), .A2(crash_dump_o_121_), .ZN(n21573) );
OR2_X1 U26383 ( .A1(n21570), .A2(crash_dump_o_119_), .ZN(n21566) );
OR2_X1 U26384 ( .A1(n21556), .A2(crash_dump_o_115_), .ZN(n21550) );
OR2_X1 U26385 ( .A1(n21547), .A2(crash_dump_o_113_), .ZN(n21543) );
OR2_X1 U26386 ( .A1(n21591), .A2(crash_dump_o_125_), .ZN(n21587) );
OR2_X1 U26387 ( .A1(n21594), .A2(crash_dump_o_126_), .ZN(n21593) );
OR2_X1 U26388 ( .A1(n21574), .A2(crash_dump_o_122_), .ZN(n21576) );
OR2_X1 U26389 ( .A1(n21567), .A2(crash_dump_o_120_), .ZN(n21569) );
OR2_X1 U26390 ( .A1(n21560), .A2(crash_dump_o_118_), .ZN(n21562) );
OR2_X1 U26391 ( .A1(n21553), .A2(crash_dump_o_116_), .ZN(n21555) );
OR2_X1 U26392 ( .A1(n21544), .A2(crash_dump_o_114_), .ZN(n21546) );
OR2_X1 U26393 ( .A1(n21537), .A2(crash_dump_o_112_), .ZN(n21539) );
OR2_X1 U26394 ( .A1(n21581), .A2(crash_dump_o_124_), .ZN(n21583) );
OR2_X1 U26395 ( .A1(n21595), .A2(crash_dump_o_127_), .ZN(n21597) );
OR2_X1 U26396 ( .A1(n6186), .A2(n11330), .ZN(n10053) );
NOR2_X1 U26397 ( .A1(n11090), .A2(n5116), .ZN(n15342) );
NAND2_X1 U26398 ( .A1(n3554), .A2(n3555), .ZN(n15737) );
OR2_X1 U26399 ( .A1(n16438), .A2(n11456), .ZN(n3554) );
NAND2_X1 U26400 ( .A1(n16437), .A2(n19962), .ZN(n3555) );
NAND2_X1 U26401 ( .A1(n7735), .A2(n7736), .ZN(n15352) );
OR2_X1 U26402 ( .A1(n16347), .A2(n11099), .ZN(n7735) );
NAND2_X1 U26403 ( .A1(n19976), .A2(n7191), .ZN(n7736) );
NOR2_X1 U26404 ( .A1(n16442), .A2(n3029), .ZN(n15739) );
NAND2_X1 U26405 ( .A1(n3030), .A2(n19884), .ZN(n3029) );
NAND2_X1 U26406 ( .A1(n11458), .A2(n3032), .ZN(n3030) );
NAND2_X1 U26407 ( .A1(n19885), .A2(n15803), .ZN(n3032) );
NOR2_X1 U26408 ( .A1(n11521), .A2(n8128), .ZN(n15783) );
NOR2_X1 U26409 ( .A1(n11292), .A2(n8128), .ZN(n15546) );
NOR2_X1 U26410 ( .A1(n11152), .A2(n8128), .ZN(n15405) );
NOR2_X1 U26411 ( .A1(n11151), .A2(n8128), .ZN(n15404) );
NOR2_X1 U26412 ( .A1(n11150), .A2(n8128), .ZN(n15403) );
NOR2_X1 U26413 ( .A1(n11149), .A2(n8128), .ZN(n15402) );
NAND2_X1 U26414 ( .A1(n2441), .A2(n2442), .ZN(n15645) );
OR2_X1 U26415 ( .A1(n1885), .A2(n11366), .ZN(n2442) );
NOR2_X1 U26416 ( .A1(n16262), .A2(n8060), .ZN(n15026) );
NOR2_X1 U26417 ( .A1(n8061), .A2(n8062), .ZN(n8060) );
NOR2_X1 U26418 ( .A1(n8056), .A2(n8063), .ZN(n8061) );
NOR2_X1 U26419 ( .A1(n10781), .A2(n16388), .ZN(n8062) );
NAND2_X1 U26420 ( .A1(n2024), .A2(n2427), .ZN(n15628) );
OR2_X1 U26421 ( .A1(n1885), .A2(n11350), .ZN(n2427) );
NAND2_X1 U26422 ( .A1(n7113), .A2(n7114), .ZN(n15182) );
OR2_X1 U26423 ( .A1(n16401), .A2(n10937), .ZN(n7114) );
NAND2_X1 U26424 ( .A1(n16400), .A2(crash_dump_o_25_), .ZN(n7113) );
NAND2_X1 U26425 ( .A1(n7123), .A2(n7124), .ZN(n15122) );
OR2_X1 U26426 ( .A1(n16401), .A2(n10877), .ZN(n7124) );
NAND2_X1 U26427 ( .A1(n16401), .A2(crash_dump_o_20_), .ZN(n7123) );
NAND2_X1 U26428 ( .A1(n7133), .A2(n7134), .ZN(n15075) );
OR2_X1 U26429 ( .A1(n16401), .A2(n10830), .ZN(n7134) );
NAND2_X1 U26430 ( .A1(n16400), .A2(crash_dump_o_16_), .ZN(n7133) );
NAND2_X1 U26431 ( .A1(crash_dump_o_66_), .A2(n19938), .ZN(n21445) );
NAND2_X1 U26432 ( .A1(n7167), .A2(n7168), .ZN(n15266) );
OR2_X1 U26433 ( .A1(n16401), .A2(n11481), .ZN(n7168) );
NAND2_X1 U26434 ( .A1(n16400), .A2(n16047), .ZN(n7167) );
NAND2_X1 U26435 ( .A1(n7170), .A2(n7171), .ZN(n15265) );
OR2_X1 U26436 ( .A1(n16401), .A2(n11487), .ZN(n7171) );
NAND2_X1 U26437 ( .A1(n16400), .A2(n16048), .ZN(n7170) );
NAND2_X1 U26438 ( .A1(n7147), .A2(n7148), .ZN(n15252) );
OR2_X1 U26439 ( .A1(n16401), .A2(n11007), .ZN(n7148) );
NAND2_X1 U26440 ( .A1(n16400), .A2(crash_dump_o_0_), .ZN(n7147) );
NAND2_X1 U26441 ( .A1(n7143), .A2(n7144), .ZN(n15223) );
OR2_X1 U26442 ( .A1(n16401), .A2(n10978), .ZN(n7144) );
NAND2_X1 U26443 ( .A1(n16400), .A2(crash_dump_o_11_), .ZN(n7143) );
NAND2_X1 U26444 ( .A1(n7109), .A2(n7110), .ZN(n15212) );
OR2_X1 U26445 ( .A1(n16401), .A2(n10967), .ZN(n7110) );
NAND2_X1 U26446 ( .A1(n16400), .A2(crash_dump_o_27_), .ZN(n7109) );
NAND2_X1 U26447 ( .A1(n7173), .A2(n7174), .ZN(n15099) );
OR2_X1 U26448 ( .A1(n16400), .A2(n10854), .ZN(n7174) );
NAND2_X1 U26449 ( .A1(n16400), .A2(n16049), .ZN(n7173) );
NAND2_X1 U26450 ( .A1(n7164), .A2(n7165), .ZN(n14920) );
OR2_X1 U26451 ( .A1(n16401), .A2(n10676), .ZN(n7165) );
NAND2_X1 U26452 ( .A1(n16400), .A2(n16050), .ZN(n7164) );
NAND2_X1 U26453 ( .A1(n7107), .A2(n7108), .ZN(n14873) );
OR2_X1 U26454 ( .A1(n16401), .A2(n10630), .ZN(n7108) );
NAND2_X1 U26455 ( .A1(n16400), .A2(crash_dump_o_28_), .ZN(n7107) );
NOR2_X1 U26456 ( .A1(n5223), .A2(n2003), .ZN(n15009) );
NOR2_X1 U26457 ( .A1(n16133), .A2(n5271), .ZN(n5223) );
NOR2_X1 U26458 ( .A1(n11310), .A2(n19970), .ZN(n15573) );
NOR2_X1 U26459 ( .A1(instr_gnt_i), .A2(n20879), .ZN(n15749) );
NAND2_X1 U26460 ( .A1(n3098), .A2(n3099), .ZN(n15725) );
OR2_X1 U26461 ( .A1(n3061), .A2(n11444), .ZN(n3099) );
NAND2_X1 U26462 ( .A1(n16438), .A2(instr_rdata_i_20_), .ZN(n3098) );
NAND2_X1 U26463 ( .A1(n3106), .A2(n3107), .ZN(n15722) );
OR2_X1 U26464 ( .A1(n16437), .A2(n11441), .ZN(n3107) );
NAND2_X1 U26465 ( .A1(n16438), .A2(instr_rdata_i_17_), .ZN(n3106) );
NAND2_X1 U26466 ( .A1(n3100), .A2(n3101), .ZN(n15706) );
OR2_X1 U26467 ( .A1(n16437), .A2(n11425), .ZN(n3101) );
NAND2_X1 U26468 ( .A1(n16438), .A2(instr_rdata_i_1_), .ZN(n3100) );
NAND2_X1 U26469 ( .A1(n2028), .A2(n2417), .ZN(n15638) );
OR2_X1 U26470 ( .A1(n1885), .A2(n11360), .ZN(n2417) );
NAND2_X1 U26471 ( .A1(n3122), .A2(n3123), .ZN(n15738) );
OR2_X1 U26472 ( .A1(n16438), .A2(n11457), .ZN(n3123) );
NAND2_X1 U26473 ( .A1(n16437), .A2(instr_rdata_i_0_), .ZN(n3122) );
NAND2_X1 U26474 ( .A1(n3074), .A2(n3075), .ZN(n15736) );
OR2_X1 U26475 ( .A1(n16438), .A2(n11455), .ZN(n3075) );
NAND2_X1 U26476 ( .A1(n3061), .A2(instr_rdata_i_31_), .ZN(n3074) );
NAND2_X1 U26477 ( .A1(n3076), .A2(n3077), .ZN(n15735) );
OR2_X1 U26478 ( .A1(n16438), .A2(n11454), .ZN(n3077) );
NAND2_X1 U26479 ( .A1(n16438), .A2(instr_rdata_i_30_), .ZN(n3076) );
NAND2_X1 U26480 ( .A1(n3080), .A2(n3081), .ZN(n15734) );
OR2_X1 U26481 ( .A1(n3061), .A2(n11453), .ZN(n3081) );
NAND2_X1 U26482 ( .A1(n3061), .A2(instr_rdata_i_29_), .ZN(n3080) );
NAND2_X1 U26483 ( .A1(n3082), .A2(n3083), .ZN(n15733) );
OR2_X1 U26484 ( .A1(n16437), .A2(n11452), .ZN(n3083) );
NAND2_X1 U26485 ( .A1(n3061), .A2(instr_rdata_i_28_), .ZN(n3082) );
NAND2_X1 U26486 ( .A1(n3084), .A2(n3085), .ZN(n15732) );
OR2_X1 U26487 ( .A1(n16437), .A2(n11451), .ZN(n3085) );
NAND2_X1 U26488 ( .A1(n16438), .A2(instr_rdata_i_27_), .ZN(n3084) );
NAND2_X1 U26489 ( .A1(n3086), .A2(n3087), .ZN(n15731) );
OR2_X1 U26490 ( .A1(n16438), .A2(n11450), .ZN(n3087) );
NAND2_X1 U26491 ( .A1(n16437), .A2(instr_rdata_i_26_), .ZN(n3086) );
NAND2_X1 U26492 ( .A1(n3088), .A2(n3089), .ZN(n15730) );
OR2_X1 U26493 ( .A1(n16438), .A2(n11449), .ZN(n3089) );
NAND2_X1 U26494 ( .A1(n16437), .A2(instr_rdata_i_25_), .ZN(n3088) );
NAND2_X1 U26495 ( .A1(n3090), .A2(n3091), .ZN(n15729) );
OR2_X1 U26496 ( .A1(n16438), .A2(n11448), .ZN(n3091) );
NAND2_X1 U26497 ( .A1(n3061), .A2(instr_rdata_i_24_), .ZN(n3090) );
NAND2_X1 U26498 ( .A1(n3092), .A2(n3093), .ZN(n15728) );
OR2_X1 U26499 ( .A1(n3061), .A2(n11447), .ZN(n3093) );
NAND2_X1 U26500 ( .A1(n16437), .A2(instr_rdata_i_23_), .ZN(n3092) );
NAND2_X1 U26501 ( .A1(n3094), .A2(n3095), .ZN(n15727) );
OR2_X1 U26502 ( .A1(n16438), .A2(n11446), .ZN(n3095) );
NAND2_X1 U26503 ( .A1(n16437), .A2(instr_rdata_i_22_), .ZN(n3094) );
NAND2_X1 U26504 ( .A1(n3096), .A2(n3097), .ZN(n15726) );
OR2_X1 U26505 ( .A1(n3061), .A2(n11445), .ZN(n3097) );
NAND2_X1 U26506 ( .A1(n16438), .A2(instr_rdata_i_21_), .ZN(n3096) );
NAND2_X1 U26507 ( .A1(n3102), .A2(n3103), .ZN(n15724) );
OR2_X1 U26508 ( .A1(n3061), .A2(n11443), .ZN(n3103) );
NAND2_X1 U26509 ( .A1(n16437), .A2(instr_rdata_i_19_), .ZN(n3102) );
NAND2_X1 U26510 ( .A1(n3104), .A2(n3105), .ZN(n15723) );
OR2_X1 U26511 ( .A1(n16437), .A2(n11442), .ZN(n3105) );
NAND2_X1 U26512 ( .A1(n16437), .A2(instr_rdata_i_18_), .ZN(n3104) );
NAND2_X1 U26513 ( .A1(n3108), .A2(n3109), .ZN(n15721) );
OR2_X1 U26514 ( .A1(n3061), .A2(n11440), .ZN(n3109) );
NAND2_X1 U26515 ( .A1(n16437), .A2(instr_rdata_i_16_), .ZN(n3108) );
NAND2_X1 U26516 ( .A1(n3110), .A2(n3111), .ZN(n15720) );
OR2_X1 U26517 ( .A1(n3061), .A2(n11439), .ZN(n3111) );
NAND2_X1 U26518 ( .A1(n16437), .A2(instr_rdata_i_15_), .ZN(n3110) );
NAND2_X1 U26519 ( .A1(n3112), .A2(n3113), .ZN(n15719) );
OR2_X1 U26520 ( .A1(n16438), .A2(n11438), .ZN(n3113) );
NAND2_X1 U26521 ( .A1(n3061), .A2(instr_rdata_i_14_), .ZN(n3112) );
NAND2_X1 U26522 ( .A1(n3114), .A2(n3115), .ZN(n15718) );
OR2_X1 U26523 ( .A1(n16437), .A2(n11437), .ZN(n3115) );
NAND2_X1 U26524 ( .A1(n16438), .A2(instr_rdata_i_13_), .ZN(n3114) );
NAND2_X1 U26525 ( .A1(n3116), .A2(n3117), .ZN(n15717) );
OR2_X1 U26526 ( .A1(n16438), .A2(n11436), .ZN(n3117) );
NAND2_X1 U26527 ( .A1(n16437), .A2(instr_rdata_i_12_), .ZN(n3116) );
NAND2_X1 U26528 ( .A1(n3118), .A2(n3119), .ZN(n15716) );
OR2_X1 U26529 ( .A1(n16438), .A2(n11435), .ZN(n3119) );
NAND2_X1 U26530 ( .A1(n3061), .A2(instr_rdata_i_11_), .ZN(n3118) );
NAND2_X1 U26531 ( .A1(n3120), .A2(n3121), .ZN(n15715) );
OR2_X1 U26532 ( .A1(n16437), .A2(n11434), .ZN(n3121) );
NAND2_X1 U26533 ( .A1(n16438), .A2(instr_rdata_i_10_), .ZN(n3120) );
NAND2_X1 U26534 ( .A1(n3059), .A2(n3060), .ZN(n15714) );
OR2_X1 U26535 ( .A1(n3061), .A2(n11433), .ZN(n3060) );
NAND2_X1 U26536 ( .A1(n3061), .A2(instr_rdata_i_9_), .ZN(n3059) );
NAND2_X1 U26537 ( .A1(n3062), .A2(n3063), .ZN(n15713) );
OR2_X1 U26538 ( .A1(n16438), .A2(n11432), .ZN(n3063) );
NAND2_X1 U26539 ( .A1(n3061), .A2(instr_rdata_i_8_), .ZN(n3062) );
NAND2_X1 U26540 ( .A1(n3064), .A2(n3065), .ZN(n15712) );
OR2_X1 U26541 ( .A1(n3061), .A2(n11431), .ZN(n3065) );
NAND2_X1 U26542 ( .A1(n16438), .A2(instr_rdata_i_7_), .ZN(n3064) );
NAND2_X1 U26543 ( .A1(n3066), .A2(n3067), .ZN(n15711) );
OR2_X1 U26544 ( .A1(n3061), .A2(n11430), .ZN(n3067) );
NAND2_X1 U26545 ( .A1(n16437), .A2(instr_rdata_i_6_), .ZN(n3066) );
NAND2_X1 U26546 ( .A1(n3068), .A2(n3069), .ZN(n15710) );
OR2_X1 U26547 ( .A1(n16437), .A2(n11429), .ZN(n3069) );
NAND2_X1 U26548 ( .A1(n16437), .A2(instr_rdata_i_5_), .ZN(n3068) );
NAND2_X1 U26549 ( .A1(n3070), .A2(n3071), .ZN(n15709) );
OR2_X1 U26550 ( .A1(n3061), .A2(n11428), .ZN(n3071) );
NAND2_X1 U26551 ( .A1(n3061), .A2(instr_rdata_i_4_), .ZN(n3070) );
NAND2_X1 U26552 ( .A1(n3072), .A2(n3073), .ZN(n15708) );
OR2_X1 U26553 ( .A1(n3061), .A2(n11427), .ZN(n3073) );
NAND2_X1 U26554 ( .A1(n16438), .A2(instr_rdata_i_3_), .ZN(n3072) );
NAND2_X1 U26555 ( .A1(n3078), .A2(n3079), .ZN(n15707) );
OR2_X1 U26556 ( .A1(n16438), .A2(n11426), .ZN(n3079) );
NAND2_X1 U26557 ( .A1(n16437), .A2(instr_rdata_i_2_), .ZN(n3078) );
NAND2_X1 U26558 ( .A1(n7767), .A2(n7768), .ZN(n15355) );
OR2_X1 U26559 ( .A1(n16347), .A2(n11102), .ZN(n7768) );
NAND2_X1 U26560 ( .A1(n19976), .A2(n7226), .ZN(n7767) );
NAND2_X1 U26561 ( .A1(n7745), .A2(n7746), .ZN(n15354) );
OR2_X1 U26562 ( .A1(n16347), .A2(n11101), .ZN(n7746) );
NAND2_X1 U26563 ( .A1(n16347), .A2(n7203), .ZN(n7745) );
NAND2_X1 U26564 ( .A1(n7739), .A2(n7740), .ZN(n15353) );
OR2_X1 U26565 ( .A1(n19976), .A2(n11100), .ZN(n7740) );
NAND2_X1 U26566 ( .A1(n19976), .A2(n7037), .ZN(n7739) );
NAND2_X1 U26567 ( .A1(n7788), .A2(n7789), .ZN(n15351) );
OR2_X1 U26568 ( .A1(n19976), .A2(n11098), .ZN(n7789) );
NAND2_X1 U26569 ( .A1(n16347), .A2(n7069), .ZN(n7788) );
NAND2_X1 U26570 ( .A1(n7786), .A2(n7787), .ZN(n15350) );
OR2_X1 U26571 ( .A1(n19976), .A2(n11097), .ZN(n7787) );
NAND2_X1 U26572 ( .A1(n19976), .A2(n7068), .ZN(n7786) );
NAND2_X1 U26573 ( .A1(n7763), .A2(n7764), .ZN(n15349) );
OR2_X1 U26574 ( .A1(n16347), .A2(n11096), .ZN(n7764) );
NAND2_X1 U26575 ( .A1(n19976), .A2(n6896), .ZN(n7763) );
NAND2_X1 U26576 ( .A1(n7741), .A2(n7742), .ZN(n15346) );
OR2_X1 U26577 ( .A1(n16347), .A2(n11093), .ZN(n7742) );
NAND2_X1 U26578 ( .A1(n19976), .A2(n6792), .ZN(n7741) );
NAND2_X1 U26579 ( .A1(n7793), .A2(n7794), .ZN(n15345) );
OR2_X1 U26580 ( .A1(n16347), .A2(n11092), .ZN(n7794) );
NAND2_X1 U26581 ( .A1(n16347), .A2(n7253), .ZN(n7793) );
NAND2_X1 U26582 ( .A1(n7751), .A2(n7752), .ZN(n15218) );
OR2_X1 U26583 ( .A1(n16347), .A2(n10973), .ZN(n7752) );
NAND2_X1 U26584 ( .A1(n19976), .A2(n6842), .ZN(n7751) );
NAND2_X1 U26585 ( .A1(n7753), .A2(n7754), .ZN(n15203) );
OR2_X1 U26586 ( .A1(n19976), .A2(n10958), .ZN(n7754) );
NAND2_X1 U26587 ( .A1(n16347), .A2(n6851), .ZN(n7753) );
NAND2_X1 U26588 ( .A1(n7755), .A2(n7756), .ZN(n15188) );
OR2_X1 U26589 ( .A1(n16347), .A2(n10943), .ZN(n7756) );
NAND2_X1 U26590 ( .A1(n16347), .A2(n6860), .ZN(n7755) );
NAND2_X1 U26591 ( .A1(n7757), .A2(n7758), .ZN(n15173) );
OR2_X1 U26592 ( .A1(n19976), .A2(n10928), .ZN(n7758) );
NAND2_X1 U26593 ( .A1(n19976), .A2(n6869), .ZN(n7757) );
NAND2_X1 U26594 ( .A1(n7759), .A2(n7760), .ZN(n15158) );
OR2_X1 U26595 ( .A1(n16347), .A2(n10913), .ZN(n7760) );
NAND2_X1 U26596 ( .A1(n16347), .A2(n6878), .ZN(n7759) );
NAND2_X1 U26597 ( .A1(n7761), .A2(n7762), .ZN(n15143) );
OR2_X1 U26598 ( .A1(n19976), .A2(n10898), .ZN(n7762) );
NAND2_X1 U26599 ( .A1(n16347), .A2(n6887), .ZN(n7761) );
NAND2_X1 U26600 ( .A1(n7765), .A2(n7766), .ZN(n15128) );
OR2_X1 U26601 ( .A1(n16347), .A2(n10883), .ZN(n7766) );
NAND2_X1 U26602 ( .A1(n19976), .A2(n6905), .ZN(n7765) );
NAND2_X1 U26603 ( .A1(n7769), .A2(n7770), .ZN(n15113) );
OR2_X1 U26604 ( .A1(n19976), .A2(n10868), .ZN(n7770) );
NAND2_X1 U26605 ( .A1(n19976), .A2(n6925), .ZN(n7769) );
NAND2_X1 U26606 ( .A1(n7771), .A2(n7772), .ZN(n15096) );
OR2_X1 U26607 ( .A1(n16347), .A2(n10851), .ZN(n7772) );
NAND2_X1 U26608 ( .A1(n16347), .A2(n6934), .ZN(n7771) );
NAND2_X1 U26609 ( .A1(n7775), .A2(n7776), .ZN(n15081) );
OR2_X1 U26610 ( .A1(n19976), .A2(n10836), .ZN(n7776) );
NAND2_X1 U26611 ( .A1(n16347), .A2(n6952), .ZN(n7775) );
NAND2_X1 U26612 ( .A1(n7728), .A2(n7729), .ZN(n14971) );
OR2_X1 U26613 ( .A1(n16347), .A2(n10727), .ZN(n7729) );
NAND2_X1 U26614 ( .A1(n19976), .A2(n7182), .ZN(n7728) );
NAND2_X1 U26615 ( .A1(n7737), .A2(n7738), .ZN(n14944) );
OR2_X1 U26616 ( .A1(n16347), .A2(n10700), .ZN(n7738) );
NAND2_X1 U26617 ( .A1(n16347), .A2(n7194), .ZN(n7737) );
NAND2_X1 U26618 ( .A1(n7730), .A2(n7731), .ZN(n14932) );
OR2_X1 U26619 ( .A1(n16347), .A2(n10688), .ZN(n7731) );
NAND2_X1 U26620 ( .A1(n19976), .A2(n7185), .ZN(n7730) );
NAND2_X1 U26621 ( .A1(n7773), .A2(n7774), .ZN(n14901) );
OR2_X1 U26622 ( .A1(n19976), .A2(n10657), .ZN(n7774) );
NAND2_X1 U26623 ( .A1(n19976), .A2(n6943), .ZN(n7773) );
NAND2_X1 U26624 ( .A1(n7749), .A2(n7750), .ZN(n14883) );
OR2_X1 U26625 ( .A1(n16347), .A2(n10640), .ZN(n7750) );
NAND2_X1 U26626 ( .A1(n16347), .A2(n6833), .ZN(n7749) );
NAND2_X1 U26627 ( .A1(n3497), .A2(n3498), .ZN(n3496) );
OR2_X1 U26628 ( .A1(n20931), .A2(n11486), .ZN(n3498) );
NOR2_X1 U26629 ( .A1(n3500), .A2(n3501), .ZN(n3497) );
NOR2_X1 U26630 ( .A1(n20753), .A2(n20926), .ZN(n3500) );
OR2_X1 U26631 ( .A1(n19938), .A2(crash_dump_o_66_), .ZN(n21444) );
NAND2_X1 U26632 ( .A1(n10985), .A2(n8079), .ZN(n15230) );
NAND2_X1 U26633 ( .A1(n2447), .A2(n2448), .ZN(n15653) );
OR2_X1 U26634 ( .A1(n1885), .A2(n11374), .ZN(n2447) );
NAND2_X1 U26635 ( .A1(n5275), .A2(n5276), .ZN(n15470) );
NAND2_X1 U26636 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_9), .ZN(n5276) );
NAND2_X1 U26637 ( .A1(n16416), .A2(n16146), .ZN(n5275) );
NAND2_X1 U26638 ( .A1(n5280), .A2(n5281), .ZN(n15469) );
NAND2_X1 U26639 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_8), .ZN(n5281) );
NAND2_X1 U26640 ( .A1(n16416), .A2(n16147), .ZN(n5280) );
NAND2_X1 U26641 ( .A1(n5283), .A2(n5284), .ZN(n15468) );
NAND2_X1 U26642 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_7), .ZN(n5284) );
NAND2_X1 U26643 ( .A1(n16416), .A2(n16148), .ZN(n5283) );
NAND2_X1 U26644 ( .A1(n5286), .A2(n5287), .ZN(n15467) );
NAND2_X1 U26645 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_6), .ZN(n5287) );
NAND2_X1 U26646 ( .A1(n16416), .A2(n16149), .ZN(n5286) );
NAND2_X1 U26647 ( .A1(n5289), .A2(n5290), .ZN(n15466) );
NAND2_X1 U26648 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_5), .ZN(n5290) );
NAND2_X1 U26649 ( .A1(n16416), .A2(n16150), .ZN(n5289) );
NAND2_X1 U26650 ( .A1(n5292), .A2(n5293), .ZN(n15465) );
NAND2_X1 U26651 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_4), .ZN(n5293) );
NAND2_X1 U26652 ( .A1(n16416), .A2(n16151), .ZN(n5292) );
NAND2_X1 U26653 ( .A1(n5295), .A2(n5296), .ZN(n15464) );
NAND2_X1 U26654 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_3), .ZN(n5296) );
NAND2_X1 U26655 ( .A1(n16416), .A2(n16152), .ZN(n5295) );
NAND2_X1 U26656 ( .A1(n5298), .A2(n5299), .ZN(n15463) );
NAND2_X1 U26657 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_31), .ZN(n5299) );
NAND2_X1 U26658 ( .A1(n16416), .A2(n16153), .ZN(n5298) );
NAND2_X1 U26659 ( .A1(n21496), .A2(n21495), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_5) );
OR2_X1 U26660 ( .A1(n21497), .A2(crash_dump_o_69_), .ZN(n21496) );
NAND2_X1 U26661 ( .A1(crash_dump_o_69_), .A2(n21497), .ZN(n21495) );
NAND2_X1 U26662 ( .A1(n22194), .A2(n22193), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_31) );
OR2_X1 U26663 ( .A1(n22198), .A2(cs_registers_i_mhpmcounter_0__31_), .ZN(n22194) );
NAND2_X1 U26664 ( .A1(cs_registers_i_mhpmcounter_0__31_), .A2(n22198), .ZN(n22193) );
NAND2_X1 U26665 ( .A1(n21453), .A2(n21452), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_21) );
OR2_X1 U26666 ( .A1(n21457), .A2(crash_dump_o_85_), .ZN(n21453) );
NAND2_X1 U26667 ( .A1(crash_dump_o_85_), .A2(n21457), .ZN(n21452) );
NAND2_X1 U26668 ( .A1(n22402), .A2(n22401), .ZN(cs_registers_i_minstret_counter_i_counter_upd_29) );
OR2_X1 U26669 ( .A1(n22409), .A2(cs_registers_i_mhpmcounter_2__29_), .ZN(n22402) );
NAND2_X1 U26670 ( .A1(cs_registers_i_mhpmcounter_2__29_), .A2(n22409), .ZN(n22401) );
NAND2_X1 U26671 ( .A1(n22224), .A2(n22223), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_3) );
OR2_X1 U26672 ( .A1(n22260), .A2(cs_registers_i_mhpmcounter_0__3_), .ZN(n22224) );
NAND2_X1 U26673 ( .A1(cs_registers_i_mhpmcounter_0__3_), .A2(n22260), .ZN(n22223) );
NAND2_X1 U26674 ( .A1(n21412), .A2(n21411), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_11) );
OR2_X1 U26675 ( .A1(n21416), .A2(crash_dump_o_75_), .ZN(n21412) );
NAND2_X1 U26676 ( .A1(crash_dump_o_75_), .A2(n21416), .ZN(n21411) );
NAND2_X1 U26677 ( .A1(n22518), .A2(n22517), .ZN(cs_registers_i_minstret_counter_i_counter_upd_5) );
OR2_X1 U26678 ( .A1(n22533), .A2(cs_registers_i_mhpmcounter_2__5_), .ZN(n22518) );
NAND2_X1 U26679 ( .A1(cs_registers_i_mhpmcounter_2__5_), .A2(n22533), .ZN(n22517) );
NAND2_X1 U26680 ( .A1(n22495), .A2(n22494), .ZN(cs_registers_i_minstret_counter_i_counter_upd_53) );
OR2_X1 U26681 ( .A1(n22499), .A2(cs_registers_i_mhpmcounter_2__53_), .ZN(n22495) );
NAND2_X1 U26682 ( .A1(cs_registers_i_mhpmcounter_2__53_), .A2(n22499), .ZN(n22494) );
NAND2_X1 U26683 ( .A1(n22433), .A2(n22432), .ZN(cs_registers_i_minstret_counter_i_counter_upd_37) );
OR2_X1 U26684 ( .A1(n22437), .A2(cs_registers_i_mhpmcounter_2__37_), .ZN(n22433) );
NAND2_X1 U26685 ( .A1(cs_registers_i_mhpmcounter_2__37_), .A2(n22437), .ZN(n22432) );
NAND2_X1 U26686 ( .A1(n22419), .A2(n22418), .ZN(cs_registers_i_minstret_counter_i_counter_upd_33) );
OR2_X1 U26687 ( .A1(n22423), .A2(cs_registers_i_mhpmcounter_2__33_), .ZN(n22419) );
NAND2_X1 U26688 ( .A1(cs_registers_i_mhpmcounter_2__33_), .A2(n22423), .ZN(n22418) );
NAND2_X1 U26689 ( .A1(n22412), .A2(n22411), .ZN(cs_registers_i_minstret_counter_i_counter_upd_31) );
OR2_X1 U26690 ( .A1(n22416), .A2(cs_registers_i_mhpmcounter_2__31_), .ZN(n22412) );
NAND2_X1 U26691 ( .A1(cs_registers_i_mhpmcounter_2__31_), .A2(n22416), .ZN(n22411) );
NAND2_X1 U26692 ( .A1(n22374), .A2(n22373), .ZN(cs_registers_i_minstret_counter_i_counter_upd_21) );
OR2_X1 U26693 ( .A1(n22378), .A2(cs_registers_i_mhpmcounter_2__21_), .ZN(n22374) );
NAND2_X1 U26694 ( .A1(cs_registers_i_mhpmcounter_2__21_), .A2(n22378), .ZN(n22373) );
NAND2_X1 U26695 ( .A1(n22300), .A2(n22299), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_5) );
OR2_X1 U26696 ( .A1(n22315), .A2(cs_registers_i_mhpmcounter_0__5_), .ZN(n22300) );
NAND2_X1 U26697 ( .A1(cs_registers_i_mhpmcounter_0__5_), .A2(n22315), .ZN(n22299) );
NAND2_X1 U26698 ( .A1(n22277), .A2(n22276), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_53) );
OR2_X1 U26699 ( .A1(n22281), .A2(cs_registers_i_mhpmcounter_0__53_), .ZN(n22277) );
NAND2_X1 U26700 ( .A1(cs_registers_i_mhpmcounter_0__53_), .A2(n22281), .ZN(n22276) );
NAND2_X1 U26701 ( .A1(n22215), .A2(n22214), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_37) );
OR2_X1 U26702 ( .A1(n22219), .A2(cs_registers_i_mhpmcounter_0__37_), .ZN(n22215) );
NAND2_X1 U26703 ( .A1(cs_registers_i_mhpmcounter_0__37_), .A2(n22219), .ZN(n22214) );
NAND2_X1 U26704 ( .A1(n22201), .A2(n22200), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_33) );
OR2_X1 U26705 ( .A1(n22205), .A2(cs_registers_i_mhpmcounter_0__33_), .ZN(n22201) );
NAND2_X1 U26706 ( .A1(cs_registers_i_mhpmcounter_0__33_), .A2(n22205), .ZN(n22200) );
NAND2_X1 U26707 ( .A1(n22156), .A2(n22155), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_21) );
OR2_X1 U26708 ( .A1(n22160), .A2(cs_registers_i_mhpmcounter_0__21_), .ZN(n22156) );
NAND2_X1 U26709 ( .A1(cs_registers_i_mhpmcounter_0__21_), .A2(n22160), .ZN(n22155) );
NAND2_X1 U26710 ( .A1(n21474), .A2(n21473), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_27) );
OR2_X1 U26711 ( .A1(n21478), .A2(crash_dump_o_91_), .ZN(n21474) );
NAND2_X1 U26712 ( .A1(crash_dump_o_91_), .A2(n21478), .ZN(n21473) );
NAND2_X1 U26713 ( .A1(n22516), .A2(n22515), .ZN(cs_registers_i_minstret_counter_i_counter_upd_59) );
OR2_X1 U26714 ( .A1(n22522), .A2(cs_registers_i_mhpmcounter_2__59_), .ZN(n22516) );
NAND2_X1 U26715 ( .A1(cs_registers_i_mhpmcounter_2__59_), .A2(n22522), .ZN(n22515) );
NAND2_X1 U26716 ( .A1(n22395), .A2(n22394), .ZN(cs_registers_i_minstret_counter_i_counter_upd_27) );
OR2_X1 U26717 ( .A1(n22399), .A2(cs_registers_i_mhpmcounter_2__27_), .ZN(n22395) );
NAND2_X1 U26718 ( .A1(cs_registers_i_mhpmcounter_2__27_), .A2(n22399), .ZN(n22394) );
NAND2_X1 U26719 ( .A1(n22298), .A2(n22297), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_59) );
OR2_X1 U26720 ( .A1(n22304), .A2(cs_registers_i_mhpmcounter_0__59_), .ZN(n22298) );
NAND2_X1 U26721 ( .A1(cs_registers_i_mhpmcounter_0__59_), .A2(n22304), .ZN(n22297) );
NAND2_X1 U26722 ( .A1(n22177), .A2(n22176), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_27) );
OR2_X1 U26723 ( .A1(n22181), .A2(cs_registers_i_mhpmcounter_0__27_), .ZN(n22177) );
NAND2_X1 U26724 ( .A1(cs_registers_i_mhpmcounter_0__27_), .A2(n22181), .ZN(n22176) );
NAND2_X1 U26725 ( .A1(n21467), .A2(n21466), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_25) );
OR2_X1 U26726 ( .A1(n21471), .A2(crash_dump_o_89_), .ZN(n21467) );
NAND2_X1 U26727 ( .A1(crash_dump_o_89_), .A2(n21471), .ZN(n21466) );
NAND2_X1 U26728 ( .A1(n22509), .A2(n22508), .ZN(cs_registers_i_minstret_counter_i_counter_upd_57) );
OR2_X1 U26729 ( .A1(n22513), .A2(cs_registers_i_mhpmcounter_2__57_), .ZN(n22509) );
NAND2_X1 U26730 ( .A1(cs_registers_i_mhpmcounter_2__57_), .A2(n22513), .ZN(n22508) );
NAND2_X1 U26731 ( .A1(n22388), .A2(n22387), .ZN(cs_registers_i_minstret_counter_i_counter_upd_25) );
OR2_X1 U26732 ( .A1(n22392), .A2(cs_registers_i_mhpmcounter_2__25_), .ZN(n22388) );
NAND2_X1 U26733 ( .A1(cs_registers_i_mhpmcounter_2__25_), .A2(n22392), .ZN(n22387) );
NAND2_X1 U26734 ( .A1(n22291), .A2(n22290), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_57) );
OR2_X1 U26735 ( .A1(n22295), .A2(cs_registers_i_mhpmcounter_0__57_), .ZN(n22291) );
NAND2_X1 U26736 ( .A1(cs_registers_i_mhpmcounter_0__57_), .A2(n22295), .ZN(n22290) );
NAND2_X1 U26737 ( .A1(n22170), .A2(n22169), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_25) );
OR2_X1 U26738 ( .A1(n22174), .A2(cs_registers_i_mhpmcounter_0__25_), .ZN(n22170) );
NAND2_X1 U26739 ( .A1(cs_registers_i_mhpmcounter_0__25_), .A2(n22174), .ZN(n22169) );
NAND2_X1 U26740 ( .A1(n21460), .A2(n21459), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_23) );
OR2_X1 U26741 ( .A1(n21464), .A2(crash_dump_o_87_), .ZN(n21460) );
NAND2_X1 U26742 ( .A1(crash_dump_o_87_), .A2(n21464), .ZN(n21459) );
NAND2_X1 U26743 ( .A1(n22502), .A2(n22501), .ZN(cs_registers_i_minstret_counter_i_counter_upd_55) );
OR2_X1 U26744 ( .A1(n22506), .A2(cs_registers_i_mhpmcounter_2__55_), .ZN(n22502) );
NAND2_X1 U26745 ( .A1(cs_registers_i_mhpmcounter_2__55_), .A2(n22506), .ZN(n22501) );
NAND2_X1 U26746 ( .A1(n22381), .A2(n22380), .ZN(cs_registers_i_minstret_counter_i_counter_upd_23) );
OR2_X1 U26747 ( .A1(n22385), .A2(cs_registers_i_mhpmcounter_2__23_), .ZN(n22381) );
NAND2_X1 U26748 ( .A1(cs_registers_i_mhpmcounter_2__23_), .A2(n22385), .ZN(n22380) );
NAND2_X1 U26749 ( .A1(n22284), .A2(n22283), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_55) );
OR2_X1 U26750 ( .A1(n22288), .A2(cs_registers_i_mhpmcounter_0__55_), .ZN(n22284) );
NAND2_X1 U26751 ( .A1(cs_registers_i_mhpmcounter_0__55_), .A2(n22288), .ZN(n22283) );
NAND2_X1 U26752 ( .A1(n22163), .A2(n22162), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_23) );
OR2_X1 U26753 ( .A1(n22167), .A2(cs_registers_i_mhpmcounter_0__23_), .ZN(n22163) );
NAND2_X1 U26754 ( .A1(cs_registers_i_mhpmcounter_0__23_), .A2(n22167), .ZN(n22162) );
NAND2_X1 U26755 ( .A1(n21440), .A2(n21439), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_19) );
OR2_X1 U26756 ( .A1(n21450), .A2(crash_dump_o_83_), .ZN(n21440) );
NAND2_X1 U26757 ( .A1(crash_dump_o_83_), .A2(n21450), .ZN(n21439) );
NAND2_X1 U26758 ( .A1(n22488), .A2(n22487), .ZN(cs_registers_i_minstret_counter_i_counter_upd_51) );
OR2_X1 U26759 ( .A1(n22492), .A2(cs_registers_i_mhpmcounter_2__51_), .ZN(n22488) );
NAND2_X1 U26760 ( .A1(cs_registers_i_mhpmcounter_2__51_), .A2(n22492), .ZN(n22487) );
NAND2_X1 U26761 ( .A1(n22365), .A2(n22364), .ZN(cs_registers_i_minstret_counter_i_counter_upd_19) );
OR2_X1 U26762 ( .A1(n22371), .A2(cs_registers_i_mhpmcounter_2__19_), .ZN(n22365) );
NAND2_X1 U26763 ( .A1(cs_registers_i_mhpmcounter_2__19_), .A2(n22371), .ZN(n22364) );
NAND2_X1 U26764 ( .A1(n22270), .A2(n22269), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_51) );
OR2_X1 U26765 ( .A1(n22274), .A2(cs_registers_i_mhpmcounter_0__51_), .ZN(n22270) );
NAND2_X1 U26766 ( .A1(cs_registers_i_mhpmcounter_0__51_), .A2(n22274), .ZN(n22269) );
NAND2_X1 U26767 ( .A1(n22147), .A2(n22146), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_19) );
OR2_X1 U26768 ( .A1(n22153), .A2(cs_registers_i_mhpmcounter_0__19_), .ZN(n22147) );
NAND2_X1 U26769 ( .A1(cs_registers_i_mhpmcounter_0__19_), .A2(n22153), .ZN(n22146) );
NAND2_X1 U26770 ( .A1(n21426), .A2(n21425), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_15) );
OR2_X1 U26771 ( .A1(n21430), .A2(crash_dump_o_79_), .ZN(n21426) );
NAND2_X1 U26772 ( .A1(crash_dump_o_79_), .A2(n21430), .ZN(n21425) );
NAND2_X1 U26773 ( .A1(n22470), .A2(n22469), .ZN(cs_registers_i_minstret_counter_i_counter_upd_47) );
OR2_X1 U26774 ( .A1(n22474), .A2(cs_registers_i_mhpmcounter_2__47_), .ZN(n22470) );
NAND2_X1 U26775 ( .A1(cs_registers_i_mhpmcounter_2__47_), .A2(n22474), .ZN(n22469) );
NAND2_X1 U26776 ( .A1(n22351), .A2(n22350), .ZN(cs_registers_i_minstret_counter_i_counter_upd_15) );
OR2_X1 U26777 ( .A1(n22355), .A2(cs_registers_i_mhpmcounter_2__15_), .ZN(n22351) );
NAND2_X1 U26778 ( .A1(cs_registers_i_mhpmcounter_2__15_), .A2(n22355), .ZN(n22350) );
NAND2_X1 U26779 ( .A1(n22252), .A2(n22251), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_47) );
OR2_X1 U26780 ( .A1(n22256), .A2(cs_registers_i_mhpmcounter_0__47_), .ZN(n22252) );
NAND2_X1 U26781 ( .A1(cs_registers_i_mhpmcounter_0__47_), .A2(n22256), .ZN(n22251) );
NAND2_X1 U26782 ( .A1(n22133), .A2(n22132), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_15) );
OR2_X1 U26783 ( .A1(n22137), .A2(cs_registers_i_mhpmcounter_0__15_), .ZN(n22133) );
NAND2_X1 U26784 ( .A1(cs_registers_i_mhpmcounter_0__15_), .A2(n22137), .ZN(n22132) );
NAND2_X1 U26785 ( .A1(n21419), .A2(n21418), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_13) );
OR2_X1 U26786 ( .A1(n21423), .A2(crash_dump_o_77_), .ZN(n21419) );
NAND2_X1 U26787 ( .A1(crash_dump_o_77_), .A2(n21423), .ZN(n21418) );
NAND2_X1 U26788 ( .A1(n22463), .A2(n22462), .ZN(cs_registers_i_minstret_counter_i_counter_upd_45) );
OR2_X1 U26789 ( .A1(n22467), .A2(cs_registers_i_mhpmcounter_2__45_), .ZN(n22463) );
NAND2_X1 U26790 ( .A1(cs_registers_i_mhpmcounter_2__45_), .A2(n22467), .ZN(n22462) );
NAND2_X1 U26791 ( .A1(n22344), .A2(n22343), .ZN(cs_registers_i_minstret_counter_i_counter_upd_13) );
OR2_X1 U26792 ( .A1(n22348), .A2(cs_registers_i_mhpmcounter_2__13_), .ZN(n22344) );
NAND2_X1 U26793 ( .A1(cs_registers_i_mhpmcounter_2__13_), .A2(n22348), .ZN(n22343) );
NAND2_X1 U26794 ( .A1(n22245), .A2(n22244), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_45) );
OR2_X1 U26795 ( .A1(n22249), .A2(cs_registers_i_mhpmcounter_0__45_), .ZN(n22245) );
NAND2_X1 U26796 ( .A1(cs_registers_i_mhpmcounter_0__45_), .A2(n22249), .ZN(n22244) );
NAND2_X1 U26797 ( .A1(n22126), .A2(n22125), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_13) );
OR2_X1 U26798 ( .A1(n22130), .A2(cs_registers_i_mhpmcounter_0__13_), .ZN(n22126) );
NAND2_X1 U26799 ( .A1(cs_registers_i_mhpmcounter_0__13_), .A2(n22130), .ZN(n22125) );
NAND2_X1 U26800 ( .A1(n22456), .A2(n22455), .ZN(cs_registers_i_minstret_counter_i_counter_upd_43) );
OR2_X1 U26801 ( .A1(n22460), .A2(cs_registers_i_mhpmcounter_2__43_), .ZN(n22456) );
NAND2_X1 U26802 ( .A1(cs_registers_i_mhpmcounter_2__43_), .A2(n22460), .ZN(n22455) );
NAND2_X1 U26803 ( .A1(n22337), .A2(n22336), .ZN(cs_registers_i_minstret_counter_i_counter_upd_11) );
OR2_X1 U26804 ( .A1(n22341), .A2(cs_registers_i_mhpmcounter_2__11_), .ZN(n22337) );
NAND2_X1 U26805 ( .A1(cs_registers_i_mhpmcounter_2__11_), .A2(n22341), .ZN(n22336) );
NAND2_X1 U26806 ( .A1(n22238), .A2(n22237), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_43) );
OR2_X1 U26807 ( .A1(n22242), .A2(cs_registers_i_mhpmcounter_0__43_), .ZN(n22238) );
NAND2_X1 U26808 ( .A1(cs_registers_i_mhpmcounter_0__43_), .A2(n22242), .ZN(n22237) );
NAND2_X1 U26809 ( .A1(n22119), .A2(n22118), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_11) );
OR2_X1 U26810 ( .A1(n22123), .A2(cs_registers_i_mhpmcounter_0__11_), .ZN(n22119) );
NAND2_X1 U26811 ( .A1(cs_registers_i_mhpmcounter_0__11_), .A2(n22123), .ZN(n22118) );
NAND2_X1 U26812 ( .A1(n21508), .A2(n21507), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_9) );
OR2_X1 U26813 ( .A1(n21509), .A2(crash_dump_o_73_), .ZN(n21508) );
NAND2_X1 U26814 ( .A1(crash_dump_o_73_), .A2(n21509), .ZN(n21507) );
NAND2_X1 U26815 ( .A1(n22449), .A2(n22448), .ZN(cs_registers_i_minstret_counter_i_counter_upd_41) );
OR2_X1 U26816 ( .A1(n22453), .A2(cs_registers_i_mhpmcounter_2__41_), .ZN(n22449) );
NAND2_X1 U26817 ( .A1(cs_registers_i_mhpmcounter_2__41_), .A2(n22453), .ZN(n22448) );
NAND2_X1 U26818 ( .A1(n22231), .A2(n22230), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_41) );
OR2_X1 U26819 ( .A1(n22235), .A2(cs_registers_i_mhpmcounter_0__41_), .ZN(n22231) );
NAND2_X1 U26820 ( .A1(cs_registers_i_mhpmcounter_0__41_), .A2(n22235), .ZN(n22230) );
NAND2_X1 U26821 ( .A1(n22538), .A2(n22537), .ZN(cs_registers_i_minstret_counter_i_counter_upd_7) );
OR2_X1 U26822 ( .A1(n22539), .A2(cs_registers_i_mhpmcounter_2__7_), .ZN(n22538) );
NAND2_X1 U26823 ( .A1(cs_registers_i_mhpmcounter_2__7_), .A2(n22539), .ZN(n22537) );
NAND2_X1 U26824 ( .A1(n22440), .A2(n22439), .ZN(cs_registers_i_minstret_counter_i_counter_upd_39) );
OR2_X1 U26825 ( .A1(n22446), .A2(cs_registers_i_mhpmcounter_2__39_), .ZN(n22440) );
NAND2_X1 U26826 ( .A1(cs_registers_i_mhpmcounter_2__39_), .A2(n22446), .ZN(n22439) );
NAND2_X1 U26827 ( .A1(n22320), .A2(n22319), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_7) );
OR2_X1 U26828 ( .A1(n22321), .A2(cs_registers_i_mhpmcounter_0__7_), .ZN(n22320) );
NAND2_X1 U26829 ( .A1(cs_registers_i_mhpmcounter_0__7_), .A2(n22321), .ZN(n22319) );
NAND2_X1 U26830 ( .A1(n22222), .A2(n22221), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_39) );
OR2_X1 U26831 ( .A1(n22228), .A2(cs_registers_i_mhpmcounter_0__39_), .ZN(n22222) );
NAND2_X1 U26832 ( .A1(cs_registers_i_mhpmcounter_0__39_), .A2(n22228), .ZN(n22221) );
NAND2_X1 U26833 ( .A1(n21502), .A2(n21501), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_7) );
OR2_X1 U26834 ( .A1(n21503), .A2(crash_dump_o_71_), .ZN(n21502) );
NAND2_X1 U26835 ( .A1(crash_dump_o_71_), .A2(n21503), .ZN(n21501) );
NAND2_X1 U26836 ( .A1(n22442), .A2(n22441), .ZN(cs_registers_i_minstret_counter_i_counter_upd_3) );
OR2_X1 U26837 ( .A1(n22478), .A2(cs_registers_i_mhpmcounter_2__3_), .ZN(n22442) );
NAND2_X1 U26838 ( .A1(cs_registers_i_mhpmcounter_2__3_), .A2(n22478), .ZN(n22441) );
NAND2_X1 U26839 ( .A1(n22426), .A2(n22425), .ZN(cs_registers_i_minstret_counter_i_counter_upd_35) );
OR2_X1 U26840 ( .A1(n22430), .A2(cs_registers_i_mhpmcounter_2__35_), .ZN(n22426) );
NAND2_X1 U26841 ( .A1(cs_registers_i_mhpmcounter_2__35_), .A2(n22430), .ZN(n22425) );
NAND2_X1 U26842 ( .A1(n22208), .A2(n22207), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_35) );
OR2_X1 U26843 ( .A1(n22212), .A2(cs_registers_i_mhpmcounter_0__35_), .ZN(n22208) );
NAND2_X1 U26844 ( .A1(cs_registers_i_mhpmcounter_0__35_), .A2(n22212), .ZN(n22207) );
NAND2_X1 U26845 ( .A1(n22477), .A2(n22476), .ZN(cs_registers_i_minstret_counter_i_counter_upd_49) );
OR2_X1 U26846 ( .A1(n22485), .A2(cs_registers_i_mhpmcounter_2__49_), .ZN(n22477) );
NAND2_X1 U26847 ( .A1(cs_registers_i_mhpmcounter_2__49_), .A2(n22485), .ZN(n22476) );
NAND2_X1 U26848 ( .A1(n22358), .A2(n22357), .ZN(cs_registers_i_minstret_counter_i_counter_upd_17) );
OR2_X1 U26849 ( .A1(n22362), .A2(cs_registers_i_mhpmcounter_2__17_), .ZN(n22358) );
NAND2_X1 U26850 ( .A1(cs_registers_i_mhpmcounter_2__17_), .A2(n22362), .ZN(n22357) );
NAND2_X1 U26851 ( .A1(n22259), .A2(n22258), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_49) );
OR2_X1 U26852 ( .A1(n22267), .A2(cs_registers_i_mhpmcounter_0__49_), .ZN(n22259) );
NAND2_X1 U26853 ( .A1(cs_registers_i_mhpmcounter_0__49_), .A2(n22267), .ZN(n22258) );
NAND2_X1 U26854 ( .A1(n22140), .A2(n22139), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_17) );
OR2_X1 U26855 ( .A1(n22144), .A2(cs_registers_i_mhpmcounter_0__17_), .ZN(n22140) );
NAND2_X1 U26856 ( .A1(cs_registers_i_mhpmcounter_0__17_), .A2(n22144), .ZN(n22139) );
NAND2_X1 U26857 ( .A1(n21433), .A2(n21432), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_17) );
OR2_X1 U26858 ( .A1(n21437), .A2(crash_dump_o_81_), .ZN(n21433) );
NAND2_X1 U26859 ( .A1(crash_dump_o_81_), .A2(n21437), .ZN(n21432) );
NAND2_X1 U26860 ( .A1(n22184), .A2(n22183), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_29) );
OR2_X1 U26861 ( .A1(n22191), .A2(cs_registers_i_mhpmcounter_0__29_), .ZN(n22184) );
NAND2_X1 U26862 ( .A1(cs_registers_i_mhpmcounter_0__29_), .A2(n22191), .ZN(n22183) );
NAND2_X1 U26863 ( .A1(n22545), .A2(n22544), .ZN(cs_registers_i_minstret_counter_i_counter_upd_9) );
OR2_X1 U26864 ( .A1(n22543), .A2(cs_registers_i_mhpmcounter_2__9_), .ZN(n22545) );
NAND2_X1 U26865 ( .A1(cs_registers_i_mhpmcounter_2__9_), .A2(n22543), .ZN(n22544) );
NAND2_X1 U26866 ( .A1(n22327), .A2(n22326), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_9) );
OR2_X1 U26867 ( .A1(n22325), .A2(cs_registers_i_mhpmcounter_0__9_), .ZN(n22327) );
NAND2_X1 U26868 ( .A1(cs_registers_i_mhpmcounter_0__9_), .A2(n22325), .ZN(n22326) );
NAND2_X1 U26869 ( .A1(n22310), .A2(n22309), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_62) );
OR2_X1 U26870 ( .A1(n22311), .A2(cs_registers_i_mhpmcounter_0__62_), .ZN(n22310) );
NAND2_X1 U26871 ( .A1(cs_registers_i_mhpmcounter_0__62_), .A2(n22311), .ZN(n22309) );
NAND2_X1 U26872 ( .A1(n21484), .A2(n21483), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_30) );
OR2_X1 U26873 ( .A1(n21487), .A2(crash_dump_o_94_), .ZN(n21484) );
NAND2_X1 U26874 ( .A1(crash_dump_o_94_), .A2(n21487), .ZN(n21483) );
NAND2_X1 U26875 ( .A1(n22525), .A2(n22524), .ZN(cs_registers_i_minstret_counter_i_counter_upd_61) );
OR2_X1 U26876 ( .A1(n22526), .A2(cs_registers_i_mhpmcounter_2__61_), .ZN(n22525) );
NAND2_X1 U26877 ( .A1(cs_registers_i_mhpmcounter_2__61_), .A2(n22526), .ZN(n22524) );
NAND2_X1 U26878 ( .A1(n22528), .A2(n22527), .ZN(cs_registers_i_minstret_counter_i_counter_upd_62) );
OR2_X1 U26879 ( .A1(n22529), .A2(cs_registers_i_mhpmcounter_2__62_), .ZN(n22528) );
NAND2_X1 U26880 ( .A1(cs_registers_i_mhpmcounter_2__62_), .A2(n22529), .ZN(n22527) );
NAND2_X1 U26881 ( .A1(n22307), .A2(n22306), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_61) );
OR2_X1 U26882 ( .A1(n22308), .A2(cs_registers_i_mhpmcounter_0__61_), .ZN(n22307) );
NAND2_X1 U26883 ( .A1(cs_registers_i_mhpmcounter_0__61_), .A2(n22308), .ZN(n22306) );
NAND2_X1 U26884 ( .A1(n21481), .A2(n21480), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_29) );
OR2_X1 U26885 ( .A1(n21482), .A2(crash_dump_o_93_), .ZN(n21481) );
NAND2_X1 U26886 ( .A1(crash_dump_o_93_), .A2(n21482), .ZN(n21480) );
NAND2_X1 U26887 ( .A1(n22367), .A2(n22366), .ZN(cs_registers_i_minstret_counter_i_counter_upd_1) );
NAND2_X1 U26888 ( .A1(cs_registers_i_mhpmcounter_2__0_), .A2(n11122), .ZN(n22367) );
NAND2_X1 U26889 ( .A1(cs_registers_i_mhpmcounter_2__1_), .A2(n11479), .ZN(n22366) );
NAND2_X1 U26890 ( .A1(n22149), .A2(n22148), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_1) );
NAND2_X1 U26891 ( .A1(cs_registers_i_mhpmcounter_0__0_), .A2(n10666), .ZN(n22149) );
NAND2_X1 U26892 ( .A1(cs_registers_i_mhpmcounter_0__1_), .A2(n10665), .ZN(n22148) );
NAND2_X1 U26893 ( .A1(n21494), .A2(n21493), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_4) );
OR2_X1 U26894 ( .A1(n21492), .A2(crash_dump_o_68_), .ZN(n21494) );
NAND2_X1 U26895 ( .A1(crash_dump_o_68_), .A2(n21492), .ZN(n21493) );
NAND2_X1 U26896 ( .A1(crash_dump_o_67_), .A2(n21491), .ZN(n21492) );
NAND2_X1 U26897 ( .A1(n21490), .A2(n21489), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_31) );
OR2_X1 U26898 ( .A1(n21488), .A2(crash_dump_o_95_), .ZN(n21490) );
NAND2_X1 U26899 ( .A1(crash_dump_o_95_), .A2(n21488), .ZN(n21489) );
NAND2_X1 U26900 ( .A1(crash_dump_o_94_), .A2(n19936), .ZN(n21488) );
NAND2_X1 U26901 ( .A1(n22532), .A2(n22531), .ZN(cs_registers_i_minstret_counter_i_counter_upd_63) );
OR2_X1 U26902 ( .A1(n22530), .A2(cs_registers_i_mhpmcounter_2__63_), .ZN(n22532) );
NAND2_X1 U26903 ( .A1(cs_registers_i_mhpmcounter_2__63_), .A2(n22530), .ZN(n22531) );
NAND2_X1 U26904 ( .A1(cs_registers_i_mhpmcounter_2__62_), .A2(n20900), .ZN(n22530) );
NAND2_X1 U26905 ( .A1(n22314), .A2(n22313), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_63) );
OR2_X1 U26906 ( .A1(n22312), .A2(cs_registers_i_mhpmcounter_0__63_), .ZN(n22314) );
NAND2_X1 U26907 ( .A1(cs_registers_i_mhpmcounter_0__63_), .A2(n22312), .ZN(n22313) );
NAND2_X1 U26908 ( .A1(cs_registers_i_mhpmcounter_0__62_), .A2(n20896), .ZN(n22312) );
NAND2_X1 U26909 ( .A1(n22405), .A2(n22404), .ZN(cs_registers_i_minstret_counter_i_counter_upd_2) );
OR2_X1 U26910 ( .A1(n22403), .A2(cs_registers_i_mhpmcounter_2__2_), .ZN(n22405) );
NAND2_X1 U26911 ( .A1(cs_registers_i_mhpmcounter_2__2_), .A2(n22403), .ZN(n22404) );
NAND2_X1 U26912 ( .A1(cs_registers_i_mhpmcounter_2__1_), .A2(cs_registers_i_mhpmcounter_2__0_), .ZN(n22403) );
NAND2_X1 U26913 ( .A1(n22187), .A2(n22186), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_2) );
OR2_X1 U26914 ( .A1(n22185), .A2(cs_registers_i_mhpmcounter_0__2_), .ZN(n22187) );
NAND2_X1 U26915 ( .A1(cs_registers_i_mhpmcounter_0__2_), .A2(n22185), .ZN(n22186) );
NAND2_X1 U26916 ( .A1(cs_registers_i_mhpmcounter_0__1_), .A2(cs_registers_i_mhpmcounter_0__0_), .ZN(n22185) );
NAND2_X1 U26917 ( .A1(n22521), .A2(n22520), .ZN(cs_registers_i_minstret_counter_i_counter_upd_60) );
OR2_X1 U26918 ( .A1(n22519), .A2(cs_registers_i_mhpmcounter_2__60_), .ZN(n22521) );
NAND2_X1 U26919 ( .A1(cs_registers_i_mhpmcounter_2__60_), .A2(n22519), .ZN(n22520) );
OR2_X1 U26920 ( .A1(n10966), .A2(n22522), .ZN(n22519) );
NAND2_X1 U26921 ( .A1(n22422), .A2(n22421), .ZN(cs_registers_i_minstret_counter_i_counter_upd_34) );
OR2_X1 U26922 ( .A1(n22420), .A2(cs_registers_i_mhpmcounter_2__34_), .ZN(n22422) );
NAND2_X1 U26923 ( .A1(cs_registers_i_mhpmcounter_2__34_), .A2(n22420), .ZN(n22421) );
OR2_X1 U26924 ( .A1(n11128), .A2(n22423), .ZN(n22420) );
NAND2_X1 U26925 ( .A1(n22415), .A2(n22414), .ZN(cs_registers_i_minstret_counter_i_counter_upd_32) );
OR2_X1 U26926 ( .A1(n22413), .A2(cs_registers_i_mhpmcounter_2__32_), .ZN(n22415) );
NAND2_X1 U26927 ( .A1(cs_registers_i_mhpmcounter_2__32_), .A2(n22413), .ZN(n22414) );
OR2_X1 U26928 ( .A1(n11126), .A2(n22416), .ZN(n22413) );
NAND2_X1 U26929 ( .A1(n22408), .A2(n22407), .ZN(cs_registers_i_minstret_counter_i_counter_upd_30) );
OR2_X1 U26930 ( .A1(n22406), .A2(cs_registers_i_mhpmcounter_2__30_), .ZN(n22408) );
NAND2_X1 U26931 ( .A1(cs_registers_i_mhpmcounter_2__30_), .A2(n22406), .ZN(n22407) );
OR2_X1 U26932 ( .A1(n11491), .A2(n22409), .ZN(n22406) );
NAND2_X1 U26933 ( .A1(n22204), .A2(n22203), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_34) );
OR2_X1 U26934 ( .A1(n22202), .A2(cs_registers_i_mhpmcounter_0__34_), .ZN(n22204) );
NAND2_X1 U26935 ( .A1(cs_registers_i_mhpmcounter_0__34_), .A2(n22202), .ZN(n22203) );
OR2_X1 U26936 ( .A1(n11117), .A2(n22205), .ZN(n22202) );
NAND2_X1 U26937 ( .A1(n22197), .A2(n22196), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_32) );
OR2_X1 U26938 ( .A1(n22195), .A2(cs_registers_i_mhpmcounter_0__32_), .ZN(n22197) );
NAND2_X1 U26939 ( .A1(cs_registers_i_mhpmcounter_0__32_), .A2(n22195), .ZN(n22196) );
OR2_X1 U26940 ( .A1(n11510), .A2(n22198), .ZN(n22195) );
NAND2_X1 U26941 ( .A1(n22190), .A2(n22189), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_30) );
OR2_X1 U26942 ( .A1(n22188), .A2(cs_registers_i_mhpmcounter_0__30_), .ZN(n22190) );
NAND2_X1 U26943 ( .A1(cs_registers_i_mhpmcounter_0__30_), .A2(n22188), .ZN(n22189) );
OR2_X1 U26944 ( .A1(n10625), .A2(n22191), .ZN(n22188) );
NAND2_X1 U26945 ( .A1(n21470), .A2(n21469), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_26) );
OR2_X1 U26946 ( .A1(n21468), .A2(crash_dump_o_90_), .ZN(n21470) );
NAND2_X1 U26947 ( .A1(crash_dump_o_90_), .A2(n21468), .ZN(n21469) );
OR2_X1 U26948 ( .A1(n10940), .A2(n21471), .ZN(n21468) );
NAND2_X1 U26949 ( .A1(n22512), .A2(n22511), .ZN(cs_registers_i_minstret_counter_i_counter_upd_58) );
OR2_X1 U26950 ( .A1(n22510), .A2(cs_registers_i_mhpmcounter_2__58_), .ZN(n22512) );
NAND2_X1 U26951 ( .A1(cs_registers_i_mhpmcounter_2__58_), .A2(n22510), .ZN(n22511) );
OR2_X1 U26952 ( .A1(n10936), .A2(n22513), .ZN(n22510) );
NAND2_X1 U26953 ( .A1(n22391), .A2(n22390), .ZN(cs_registers_i_minstret_counter_i_counter_upd_26) );
OR2_X1 U26954 ( .A1(n22389), .A2(cs_registers_i_mhpmcounter_2__26_), .ZN(n22391) );
NAND2_X1 U26955 ( .A1(cs_registers_i_mhpmcounter_2__26_), .A2(n22389), .ZN(n22390) );
OR2_X1 U26956 ( .A1(n10935), .A2(n22392), .ZN(n22389) );
NAND2_X1 U26957 ( .A1(n22294), .A2(n22293), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_58) );
OR2_X1 U26958 ( .A1(n22292), .A2(cs_registers_i_mhpmcounter_0__58_), .ZN(n22294) );
NAND2_X1 U26959 ( .A1(cs_registers_i_mhpmcounter_0__58_), .A2(n22292), .ZN(n22293) );
OR2_X1 U26960 ( .A1(n10934), .A2(n22295), .ZN(n22292) );
NAND2_X1 U26961 ( .A1(n22173), .A2(n22172), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_26) );
OR2_X1 U26962 ( .A1(n22171), .A2(cs_registers_i_mhpmcounter_0__26_), .ZN(n22173) );
NAND2_X1 U26963 ( .A1(cs_registers_i_mhpmcounter_0__26_), .A2(n22171), .ZN(n22172) );
OR2_X1 U26964 ( .A1(n10933), .A2(n22174), .ZN(n22171) );
NAND2_X1 U26965 ( .A1(n21463), .A2(n21462), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_24) );
OR2_X1 U26966 ( .A1(n21461), .A2(crash_dump_o_88_), .ZN(n21463) );
NAND2_X1 U26967 ( .A1(crash_dump_o_88_), .A2(n21461), .ZN(n21462) );
OR2_X1 U26968 ( .A1(n10910), .A2(n21464), .ZN(n21461) );
NAND2_X1 U26969 ( .A1(n22505), .A2(n22504), .ZN(cs_registers_i_minstret_counter_i_counter_upd_56) );
OR2_X1 U26970 ( .A1(n22503), .A2(cs_registers_i_mhpmcounter_2__56_), .ZN(n22505) );
NAND2_X1 U26971 ( .A1(cs_registers_i_mhpmcounter_2__56_), .A2(n22503), .ZN(n22504) );
OR2_X1 U26972 ( .A1(n10906), .A2(n22506), .ZN(n22503) );
NAND2_X1 U26973 ( .A1(n22384), .A2(n22383), .ZN(cs_registers_i_minstret_counter_i_counter_upd_24) );
OR2_X1 U26974 ( .A1(n22382), .A2(cs_registers_i_mhpmcounter_2__24_), .ZN(n22384) );
NAND2_X1 U26975 ( .A1(cs_registers_i_mhpmcounter_2__24_), .A2(n22382), .ZN(n22383) );
OR2_X1 U26976 ( .A1(n10905), .A2(n22385), .ZN(n22382) );
NAND2_X1 U26977 ( .A1(n22287), .A2(n22286), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_56) );
OR2_X1 U26978 ( .A1(n22285), .A2(cs_registers_i_mhpmcounter_0__56_), .ZN(n22287) );
NAND2_X1 U26979 ( .A1(cs_registers_i_mhpmcounter_0__56_), .A2(n22285), .ZN(n22286) );
OR2_X1 U26980 ( .A1(n10904), .A2(n22288), .ZN(n22285) );
NAND2_X1 U26981 ( .A1(n22166), .A2(n22165), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_24) );
OR2_X1 U26982 ( .A1(n22164), .A2(cs_registers_i_mhpmcounter_0__24_), .ZN(n22166) );
NAND2_X1 U26983 ( .A1(cs_registers_i_mhpmcounter_0__24_), .A2(n22164), .ZN(n22165) );
OR2_X1 U26984 ( .A1(n10903), .A2(n22167), .ZN(n22164) );
NAND2_X1 U26985 ( .A1(n21456), .A2(n21455), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_22) );
OR2_X1 U26986 ( .A1(n21454), .A2(crash_dump_o_86_), .ZN(n21456) );
NAND2_X1 U26987 ( .A1(crash_dump_o_86_), .A2(n21454), .ZN(n21455) );
OR2_X1 U26988 ( .A1(n11496), .A2(n21457), .ZN(n21454) );
NAND2_X1 U26989 ( .A1(n22498), .A2(n22497), .ZN(cs_registers_i_minstret_counter_i_counter_upd_54) );
OR2_X1 U26990 ( .A1(n22496), .A2(cs_registers_i_mhpmcounter_2__54_), .ZN(n22498) );
NAND2_X1 U26991 ( .A1(cs_registers_i_mhpmcounter_2__54_), .A2(n22496), .ZN(n22497) );
OR2_X1 U26992 ( .A1(n11131), .A2(n22499), .ZN(n22496) );
NAND2_X1 U26993 ( .A1(n22377), .A2(n22376), .ZN(cs_registers_i_minstret_counter_i_counter_upd_22) );
OR2_X1 U26994 ( .A1(n22375), .A2(cs_registers_i_mhpmcounter_2__22_), .ZN(n22377) );
NAND2_X1 U26995 ( .A1(cs_registers_i_mhpmcounter_2__22_), .A2(n22375), .ZN(n22376) );
OR2_X1 U26996 ( .A1(n11123), .A2(n22378), .ZN(n22375) );
NAND2_X1 U26997 ( .A1(n22280), .A2(n22279), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_54) );
OR2_X1 U26998 ( .A1(n22278), .A2(cs_registers_i_mhpmcounter_0__54_), .ZN(n22280) );
NAND2_X1 U26999 ( .A1(cs_registers_i_mhpmcounter_0__54_), .A2(n22278), .ZN(n22279) );
OR2_X1 U27000 ( .A1(n11120), .A2(n22281), .ZN(n22278) );
NAND2_X1 U27001 ( .A1(n22159), .A2(n22158), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_22) );
OR2_X1 U27002 ( .A1(n22157), .A2(cs_registers_i_mhpmcounter_0__22_), .ZN(n22159) );
NAND2_X1 U27003 ( .A1(cs_registers_i_mhpmcounter_0__22_), .A2(n22157), .ZN(n22158) );
OR2_X1 U27004 ( .A1(n11114), .A2(n22160), .ZN(n22157) );
NAND2_X1 U27005 ( .A1(n21443), .A2(n21442), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_20) );
OR2_X1 U27006 ( .A1(n21441), .A2(crash_dump_o_84_), .ZN(n21443) );
NAND2_X1 U27007 ( .A1(crash_dump_o_84_), .A2(n21441), .ZN(n21442) );
OR2_X1 U27008 ( .A1(n10865), .A2(n21450), .ZN(n21441) );
NAND2_X1 U27009 ( .A1(n22491), .A2(n22490), .ZN(cs_registers_i_minstret_counter_i_counter_upd_52) );
OR2_X1 U27010 ( .A1(n22489), .A2(cs_registers_i_mhpmcounter_2__52_), .ZN(n22491) );
NAND2_X1 U27011 ( .A1(cs_registers_i_mhpmcounter_2__52_), .A2(n22489), .ZN(n22490) );
OR2_X1 U27012 ( .A1(n10861), .A2(n22492), .ZN(n22489) );
NAND2_X1 U27013 ( .A1(n22370), .A2(n22369), .ZN(cs_registers_i_minstret_counter_i_counter_upd_20) );
OR2_X1 U27014 ( .A1(n22368), .A2(cs_registers_i_mhpmcounter_2__20_), .ZN(n22370) );
NAND2_X1 U27015 ( .A1(cs_registers_i_mhpmcounter_2__20_), .A2(n22368), .ZN(n22369) );
OR2_X1 U27016 ( .A1(n10860), .A2(n22371), .ZN(n22368) );
NAND2_X1 U27017 ( .A1(n22273), .A2(n22272), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_52) );
OR2_X1 U27018 ( .A1(n22271), .A2(cs_registers_i_mhpmcounter_0__52_), .ZN(n22273) );
NAND2_X1 U27019 ( .A1(cs_registers_i_mhpmcounter_0__52_), .A2(n22271), .ZN(n22272) );
OR2_X1 U27020 ( .A1(n10859), .A2(n22274), .ZN(n22271) );
NAND2_X1 U27021 ( .A1(n22152), .A2(n22151), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_20) );
OR2_X1 U27022 ( .A1(n22150), .A2(cs_registers_i_mhpmcounter_0__20_), .ZN(n22152) );
NAND2_X1 U27023 ( .A1(cs_registers_i_mhpmcounter_0__20_), .A2(n22150), .ZN(n22151) );
OR2_X1 U27024 ( .A1(n10858), .A2(n22153), .ZN(n22150) );
NAND2_X1 U27025 ( .A1(n21436), .A2(n21435), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_18) );
OR2_X1 U27026 ( .A1(n21434), .A2(crash_dump_o_82_), .ZN(n21436) );
NAND2_X1 U27027 ( .A1(crash_dump_o_82_), .A2(n21434), .ZN(n21435) );
OR2_X1 U27028 ( .A1(n10648), .A2(n21437), .ZN(n21434) );
NAND2_X1 U27029 ( .A1(n22484), .A2(n22483), .ZN(cs_registers_i_minstret_counter_i_counter_upd_50) );
OR2_X1 U27030 ( .A1(n22482), .A2(cs_registers_i_mhpmcounter_2__50_), .ZN(n22484) );
NAND2_X1 U27031 ( .A1(cs_registers_i_mhpmcounter_2__50_), .A2(n22482), .ZN(n22483) );
OR2_X1 U27032 ( .A1(n10653), .A2(n22485), .ZN(n22482) );
NAND2_X1 U27033 ( .A1(n22361), .A2(n22360), .ZN(cs_registers_i_minstret_counter_i_counter_upd_18) );
OR2_X1 U27034 ( .A1(n22359), .A2(cs_registers_i_mhpmcounter_2__18_), .ZN(n22361) );
NAND2_X1 U27035 ( .A1(cs_registers_i_mhpmcounter_2__18_), .A2(n22359), .ZN(n22360) );
OR2_X1 U27036 ( .A1(n10652), .A2(n22362), .ZN(n22359) );
NAND2_X1 U27037 ( .A1(n22266), .A2(n22265), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_50) );
OR2_X1 U27038 ( .A1(n22264), .A2(cs_registers_i_mhpmcounter_0__50_), .ZN(n22266) );
NAND2_X1 U27039 ( .A1(cs_registers_i_mhpmcounter_0__50_), .A2(n22264), .ZN(n22265) );
OR2_X1 U27040 ( .A1(n10651), .A2(n22267), .ZN(n22264) );
NAND2_X1 U27041 ( .A1(n22143), .A2(n22142), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_18) );
OR2_X1 U27042 ( .A1(n22141), .A2(cs_registers_i_mhpmcounter_0__18_), .ZN(n22143) );
NAND2_X1 U27043 ( .A1(cs_registers_i_mhpmcounter_0__18_), .A2(n22141), .ZN(n22142) );
OR2_X1 U27044 ( .A1(n10650), .A2(n22144), .ZN(n22141) );
NAND2_X1 U27045 ( .A1(n21429), .A2(n21428), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_16) );
OR2_X1 U27046 ( .A1(n21427), .A2(crash_dump_o_80_), .ZN(n21429) );
NAND2_X1 U27047 ( .A1(crash_dump_o_80_), .A2(n21427), .ZN(n21428) );
OR2_X1 U27048 ( .A1(n10818), .A2(n21430), .ZN(n21427) );
NAND2_X1 U27049 ( .A1(n22473), .A2(n22472), .ZN(cs_registers_i_minstret_counter_i_counter_upd_48) );
OR2_X1 U27050 ( .A1(n22471), .A2(cs_registers_i_mhpmcounter_2__48_), .ZN(n22473) );
NAND2_X1 U27051 ( .A1(cs_registers_i_mhpmcounter_2__48_), .A2(n22471), .ZN(n22472) );
OR2_X1 U27052 ( .A1(n10814), .A2(n22474), .ZN(n22471) );
NAND2_X1 U27053 ( .A1(n22354), .A2(n22353), .ZN(cs_registers_i_minstret_counter_i_counter_upd_16) );
OR2_X1 U27054 ( .A1(n22352), .A2(cs_registers_i_mhpmcounter_2__16_), .ZN(n22354) );
NAND2_X1 U27055 ( .A1(cs_registers_i_mhpmcounter_2__16_), .A2(n22352), .ZN(n22353) );
OR2_X1 U27056 ( .A1(n10813), .A2(n22355), .ZN(n22352) );
NAND2_X1 U27057 ( .A1(n22255), .A2(n22254), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_48) );
OR2_X1 U27058 ( .A1(n22253), .A2(cs_registers_i_mhpmcounter_0__48_), .ZN(n22255) );
NAND2_X1 U27059 ( .A1(cs_registers_i_mhpmcounter_0__48_), .A2(n22253), .ZN(n22254) );
OR2_X1 U27060 ( .A1(n10812), .A2(n22256), .ZN(n22253) );
NAND2_X1 U27061 ( .A1(n22136), .A2(n22135), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_16) );
OR2_X1 U27062 ( .A1(n22134), .A2(cs_registers_i_mhpmcounter_0__16_), .ZN(n22136) );
NAND2_X1 U27063 ( .A1(cs_registers_i_mhpmcounter_0__16_), .A2(n22134), .ZN(n22135) );
OR2_X1 U27064 ( .A1(n10811), .A2(n22137), .ZN(n22134) );
NAND2_X1 U27065 ( .A1(n21422), .A2(n21421), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_14) );
OR2_X1 U27066 ( .A1(n21420), .A2(crash_dump_o_78_), .ZN(n21422) );
NAND2_X1 U27067 ( .A1(crash_dump_o_78_), .A2(n21420), .ZN(n21421) );
OR2_X1 U27068 ( .A1(n10789), .A2(n21423), .ZN(n21420) );
NAND2_X1 U27069 ( .A1(n22466), .A2(n22465), .ZN(cs_registers_i_minstret_counter_i_counter_upd_46) );
OR2_X1 U27070 ( .A1(n22464), .A2(cs_registers_i_mhpmcounter_2__46_), .ZN(n22466) );
NAND2_X1 U27071 ( .A1(cs_registers_i_mhpmcounter_2__46_), .A2(n22464), .ZN(n22465) );
OR2_X1 U27072 ( .A1(n10785), .A2(n22467), .ZN(n22464) );
NAND2_X1 U27073 ( .A1(n22347), .A2(n22346), .ZN(cs_registers_i_minstret_counter_i_counter_upd_14) );
OR2_X1 U27074 ( .A1(n22345), .A2(cs_registers_i_mhpmcounter_2__14_), .ZN(n22347) );
NAND2_X1 U27075 ( .A1(cs_registers_i_mhpmcounter_2__14_), .A2(n22345), .ZN(n22346) );
OR2_X1 U27076 ( .A1(n10784), .A2(n22348), .ZN(n22345) );
NAND2_X1 U27077 ( .A1(n22248), .A2(n22247), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_46) );
OR2_X1 U27078 ( .A1(n22246), .A2(cs_registers_i_mhpmcounter_0__46_), .ZN(n22248) );
NAND2_X1 U27079 ( .A1(cs_registers_i_mhpmcounter_0__46_), .A2(n22246), .ZN(n22247) );
OR2_X1 U27080 ( .A1(n10783), .A2(n22249), .ZN(n22246) );
NAND2_X1 U27081 ( .A1(n22129), .A2(n22128), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_14) );
OR2_X1 U27082 ( .A1(n22127), .A2(cs_registers_i_mhpmcounter_0__14_), .ZN(n22129) );
NAND2_X1 U27083 ( .A1(cs_registers_i_mhpmcounter_0__14_), .A2(n22127), .ZN(n22128) );
OR2_X1 U27084 ( .A1(n10782), .A2(n22130), .ZN(n22127) );
NAND2_X1 U27085 ( .A1(n22459), .A2(n22458), .ZN(cs_registers_i_minstret_counter_i_counter_upd_44) );
OR2_X1 U27086 ( .A1(n22457), .A2(cs_registers_i_mhpmcounter_2__44_), .ZN(n22459) );
NAND2_X1 U27087 ( .A1(cs_registers_i_mhpmcounter_2__44_), .A2(n22457), .ZN(n22458) );
OR2_X1 U27088 ( .A1(n10764), .A2(n22460), .ZN(n22457) );
NAND2_X1 U27089 ( .A1(n22340), .A2(n22339), .ZN(cs_registers_i_minstret_counter_i_counter_upd_12) );
OR2_X1 U27090 ( .A1(n22338), .A2(cs_registers_i_mhpmcounter_2__12_), .ZN(n22340) );
NAND2_X1 U27091 ( .A1(cs_registers_i_mhpmcounter_2__12_), .A2(n22338), .ZN(n22339) );
OR2_X1 U27092 ( .A1(n10763), .A2(n22341), .ZN(n22338) );
NAND2_X1 U27093 ( .A1(n22241), .A2(n22240), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_44) );
OR2_X1 U27094 ( .A1(n22239), .A2(cs_registers_i_mhpmcounter_0__44_), .ZN(n22241) );
NAND2_X1 U27095 ( .A1(cs_registers_i_mhpmcounter_0__44_), .A2(n22239), .ZN(n22240) );
OR2_X1 U27096 ( .A1(n10762), .A2(n22242), .ZN(n22239) );
NAND2_X1 U27097 ( .A1(n22122), .A2(n22121), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_12) );
OR2_X1 U27098 ( .A1(n22120), .A2(cs_registers_i_mhpmcounter_0__12_), .ZN(n22122) );
NAND2_X1 U27099 ( .A1(cs_registers_i_mhpmcounter_0__12_), .A2(n22120), .ZN(n22121) );
OR2_X1 U27100 ( .A1(n10761), .A2(n22123), .ZN(n22120) );
NAND2_X1 U27101 ( .A1(n21415), .A2(n21414), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_12) );
OR2_X1 U27102 ( .A1(n21413), .A2(crash_dump_o_76_), .ZN(n21415) );
NAND2_X1 U27103 ( .A1(crash_dump_o_76_), .A2(n21413), .ZN(n21414) );
OR2_X1 U27104 ( .A1(n11308), .A2(n21416), .ZN(n21413) );
NAND2_X1 U27105 ( .A1(n21512), .A2(n21511), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_10) );
OR2_X1 U27106 ( .A1(n21510), .A2(crash_dump_o_74_), .ZN(n21512) );
NAND2_X1 U27107 ( .A1(crash_dump_o_74_), .A2(n21510), .ZN(n21511) );
OR2_X1 U27108 ( .A1(n10746), .A2(n21509), .ZN(n21510) );
NAND2_X1 U27109 ( .A1(n22452), .A2(n22451), .ZN(cs_registers_i_minstret_counter_i_counter_upd_42) );
OR2_X1 U27110 ( .A1(n22450), .A2(cs_registers_i_mhpmcounter_2__42_), .ZN(n22452) );
NAND2_X1 U27111 ( .A1(cs_registers_i_mhpmcounter_2__42_), .A2(n22450), .ZN(n22451) );
OR2_X1 U27112 ( .A1(n10735), .A2(n22453), .ZN(n22450) );
NAND2_X1 U27113 ( .A1(n22234), .A2(n22233), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_42) );
OR2_X1 U27114 ( .A1(n22232), .A2(cs_registers_i_mhpmcounter_0__42_), .ZN(n22234) );
NAND2_X1 U27115 ( .A1(cs_registers_i_mhpmcounter_0__42_), .A2(n22232), .ZN(n22233) );
OR2_X1 U27116 ( .A1(n10733), .A2(n22235), .ZN(n22232) );
NAND2_X1 U27117 ( .A1(n21506), .A2(n21505), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_8) );
OR2_X1 U27118 ( .A1(n21504), .A2(crash_dump_o_72_), .ZN(n21506) );
NAND2_X1 U27119 ( .A1(crash_dump_o_72_), .A2(n21504), .ZN(n21505) );
OR2_X1 U27120 ( .A1(n10681), .A2(n21503), .ZN(n21504) );
NAND2_X1 U27121 ( .A1(n22542), .A2(n22541), .ZN(cs_registers_i_minstret_counter_i_counter_upd_8) );
OR2_X1 U27122 ( .A1(n22540), .A2(cs_registers_i_mhpmcounter_2__8_), .ZN(n22542) );
NAND2_X1 U27123 ( .A1(cs_registers_i_mhpmcounter_2__8_), .A2(n22540), .ZN(n22541) );
OR2_X1 U27124 ( .A1(n10686), .A2(n22539), .ZN(n22540) );
NAND2_X1 U27125 ( .A1(n22445), .A2(n22444), .ZN(cs_registers_i_minstret_counter_i_counter_upd_40) );
OR2_X1 U27126 ( .A1(n22443), .A2(cs_registers_i_mhpmcounter_2__40_), .ZN(n22445) );
NAND2_X1 U27127 ( .A1(cs_registers_i_mhpmcounter_2__40_), .A2(n22443), .ZN(n22444) );
OR2_X1 U27128 ( .A1(n10685), .A2(n22446), .ZN(n22443) );
NAND2_X1 U27129 ( .A1(n22324), .A2(n22323), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_8) );
OR2_X1 U27130 ( .A1(n22322), .A2(cs_registers_i_mhpmcounter_0__8_), .ZN(n22324) );
NAND2_X1 U27131 ( .A1(cs_registers_i_mhpmcounter_0__8_), .A2(n22322), .ZN(n22323) );
OR2_X1 U27132 ( .A1(n10684), .A2(n22321), .ZN(n22322) );
NAND2_X1 U27133 ( .A1(n22227), .A2(n22226), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_40) );
OR2_X1 U27134 ( .A1(n22225), .A2(cs_registers_i_mhpmcounter_0__40_), .ZN(n22227) );
NAND2_X1 U27135 ( .A1(cs_registers_i_mhpmcounter_0__40_), .A2(n22225), .ZN(n22226) );
OR2_X1 U27136 ( .A1(n10683), .A2(n22228), .ZN(n22225) );
NAND2_X1 U27137 ( .A1(n21500), .A2(n21499), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_6) );
OR2_X1 U27138 ( .A1(n21498), .A2(crash_dump_o_70_), .ZN(n21500) );
NAND2_X1 U27139 ( .A1(crash_dump_o_70_), .A2(n21498), .ZN(n21499) );
OR2_X1 U27140 ( .A1(n11513), .A2(n21497), .ZN(n21498) );
NAND2_X1 U27141 ( .A1(n22536), .A2(n22535), .ZN(cs_registers_i_minstret_counter_i_counter_upd_6) );
OR2_X1 U27142 ( .A1(n22534), .A2(cs_registers_i_mhpmcounter_2__6_), .ZN(n22536) );
NAND2_X1 U27143 ( .A1(cs_registers_i_mhpmcounter_2__6_), .A2(n22534), .ZN(n22535) );
OR2_X1 U27144 ( .A1(n11132), .A2(n22533), .ZN(n22534) );
NAND2_X1 U27145 ( .A1(n22436), .A2(n22435), .ZN(cs_registers_i_minstret_counter_i_counter_upd_38) );
OR2_X1 U27146 ( .A1(n22434), .A2(cs_registers_i_mhpmcounter_2__38_), .ZN(n22436) );
NAND2_X1 U27147 ( .A1(cs_registers_i_mhpmcounter_2__38_), .A2(n22434), .ZN(n22435) );
OR2_X1 U27148 ( .A1(n11130), .A2(n22437), .ZN(n22434) );
NAND2_X1 U27149 ( .A1(n22318), .A2(n22317), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_6) );
OR2_X1 U27150 ( .A1(n22316), .A2(cs_registers_i_mhpmcounter_0__6_), .ZN(n22318) );
NAND2_X1 U27151 ( .A1(cs_registers_i_mhpmcounter_0__6_), .A2(n22316), .ZN(n22317) );
OR2_X1 U27152 ( .A1(n11121), .A2(n22315), .ZN(n22316) );
NAND2_X1 U27153 ( .A1(n22218), .A2(n22217), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_38) );
OR2_X1 U27154 ( .A1(n22216), .A2(cs_registers_i_mhpmcounter_0__38_), .ZN(n22218) );
NAND2_X1 U27155 ( .A1(cs_registers_i_mhpmcounter_0__38_), .A2(n22216), .ZN(n22217) );
OR2_X1 U27156 ( .A1(n11119), .A2(n22219), .ZN(n22216) );
NAND2_X1 U27157 ( .A1(n22481), .A2(n22480), .ZN(cs_registers_i_minstret_counter_i_counter_upd_4) );
OR2_X1 U27158 ( .A1(n22479), .A2(cs_registers_i_mhpmcounter_2__4_), .ZN(n22481) );
NAND2_X1 U27159 ( .A1(cs_registers_i_mhpmcounter_2__4_), .A2(n22479), .ZN(n22480) );
OR2_X1 U27160 ( .A1(n10675), .A2(n22478), .ZN(n22479) );
NAND2_X1 U27161 ( .A1(n22429), .A2(n22428), .ZN(cs_registers_i_minstret_counter_i_counter_upd_36) );
OR2_X1 U27162 ( .A1(n22427), .A2(cs_registers_i_mhpmcounter_2__36_), .ZN(n22429) );
NAND2_X1 U27163 ( .A1(cs_registers_i_mhpmcounter_2__36_), .A2(n22427), .ZN(n22428) );
OR2_X1 U27164 ( .A1(n10674), .A2(n22430), .ZN(n22427) );
NAND2_X1 U27165 ( .A1(n22263), .A2(n22262), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_4) );
OR2_X1 U27166 ( .A1(n22261), .A2(cs_registers_i_mhpmcounter_0__4_), .ZN(n22263) );
NAND2_X1 U27167 ( .A1(cs_registers_i_mhpmcounter_0__4_), .A2(n22261), .ZN(n22262) );
OR2_X1 U27168 ( .A1(n11478), .A2(n22260), .ZN(n22261) );
NAND2_X1 U27169 ( .A1(n22211), .A2(n22210), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_36) );
OR2_X1 U27170 ( .A1(n22209), .A2(cs_registers_i_mhpmcounter_0__36_), .ZN(n22211) );
NAND2_X1 U27171 ( .A1(cs_registers_i_mhpmcounter_0__36_), .A2(n22209), .ZN(n22210) );
OR2_X1 U27172 ( .A1(n10673), .A2(n22212), .ZN(n22209) );
NAND2_X1 U27173 ( .A1(n22398), .A2(n22397), .ZN(cs_registers_i_minstret_counter_i_counter_upd_28) );
OR2_X1 U27174 ( .A1(n22396), .A2(cs_registers_i_mhpmcounter_2__28_), .ZN(n22398) );
NAND2_X1 U27175 ( .A1(cs_registers_i_mhpmcounter_2__28_), .A2(n22396), .ZN(n22397) );
OR2_X1 U27176 ( .A1(n10965), .A2(n22399), .ZN(n22396) );
NAND2_X1 U27177 ( .A1(n22303), .A2(n22302), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_60) );
OR2_X1 U27178 ( .A1(n22301), .A2(cs_registers_i_mhpmcounter_0__60_), .ZN(n22303) );
NAND2_X1 U27179 ( .A1(cs_registers_i_mhpmcounter_0__60_), .A2(n22301), .ZN(n22302) );
OR2_X1 U27180 ( .A1(n10964), .A2(n22304), .ZN(n22301) );
NAND2_X1 U27181 ( .A1(n22180), .A2(n22179), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_28) );
OR2_X1 U27182 ( .A1(n22178), .A2(cs_registers_i_mhpmcounter_0__28_), .ZN(n22180) );
NAND2_X1 U27183 ( .A1(cs_registers_i_mhpmcounter_0__28_), .A2(n22178), .ZN(n22179) );
OR2_X1 U27184 ( .A1(n10963), .A2(n22181), .ZN(n22178) );
NAND2_X1 U27185 ( .A1(n21477), .A2(n21476), .ZN(if_stage_i_gen_prefetch_buffer_prefetch_buffer_i_addr_next_28) );
OR2_X1 U27186 ( .A1(n21475), .A2(crash_dump_o_92_), .ZN(n21477) );
NAND2_X1 U27187 ( .A1(crash_dump_o_92_), .A2(n21475), .ZN(n21476) );
OR2_X1 U27188 ( .A1(n10970), .A2(n21478), .ZN(n21475) );
NAND2_X1 U27189 ( .A1(n22334), .A2(n22333), .ZN(cs_registers_i_minstret_counter_i_counter_upd_10) );
OR2_X1 U27190 ( .A1(n22332), .A2(cs_registers_i_mhpmcounter_2__10_), .ZN(n22334) );
NAND2_X1 U27191 ( .A1(cs_registers_i_mhpmcounter_2__10_), .A2(n22332), .ZN(n22333) );
OR2_X1 U27192 ( .A1(n22543), .A2(n10736), .ZN(n22332) );
NAND2_X1 U27193 ( .A1(n22116), .A2(n22115), .ZN(cs_registers_i_mcycle_counter_i_counter_upd_10) );
OR2_X1 U27194 ( .A1(n22114), .A2(cs_registers_i_mhpmcounter_0__10_), .ZN(n22116) );
NAND2_X1 U27195 ( .A1(cs_registers_i_mhpmcounter_0__10_), .A2(n22114), .ZN(n22115) );
OR2_X1 U27196 ( .A1(n22325), .A2(n10734), .ZN(n22114) );
NAND2_X1 U27197 ( .A1(n3010), .A2(n3011), .ZN(n14832) );
NOR2_X1 U27198 ( .A1(n3012), .A2(n3013), .ZN(n3010) );
NAND2_X1 U27199 ( .A1(n16445), .A2(n16051), .ZN(n3011) );
NOR2_X1 U27200 ( .A1(n10590), .A2(n16444), .ZN(n3012) );
NAND2_X1 U27201 ( .A1(n1958), .A2(n1959), .ZN(n15744) );
OR2_X1 U27202 ( .A1(n1885), .A2(n11465), .ZN(n1958) );
NAND2_X1 U27203 ( .A1(n16452), .A2(crash_dump_o_65_), .ZN(n1959) );
NAND2_X1 U27204 ( .A1(n2445), .A2(n2446), .ZN(n15742) );
OR2_X1 U27205 ( .A1(n16450), .A2(n11463), .ZN(n2445) );
NAND2_X1 U27206 ( .A1(n16452), .A2(n2275), .ZN(n2446) );
NAND2_X1 U27207 ( .A1(n2433), .A2(n2434), .ZN(n15651) );
OR2_X1 U27208 ( .A1(n16450), .A2(n11372), .ZN(n2433) );
NAND2_X1 U27209 ( .A1(n16453), .A2(n2035), .ZN(n2434) );
NAND2_X1 U27210 ( .A1(n2435), .A2(n2436), .ZN(n15649) );
OR2_X1 U27211 ( .A1(n1885), .A2(n11370), .ZN(n2435) );
NAND2_X1 U27212 ( .A1(n16451), .A2(n2437), .ZN(n2436) );
NAND2_X1 U27213 ( .A1(n2438), .A2(n2439), .ZN(n15647) );
OR2_X1 U27214 ( .A1(n16453), .A2(n11368), .ZN(n2438) );
NAND2_X1 U27215 ( .A1(n16451), .A2(n2440), .ZN(n2439) );
NAND2_X1 U27216 ( .A1(n2443), .A2(n2444), .ZN(n15643) );
OR2_X1 U27217 ( .A1(n16453), .A2(n11364), .ZN(n2443) );
NAND2_X1 U27218 ( .A1(n16450), .A2(n2103), .ZN(n2444) );
NAND2_X1 U27219 ( .A1(n2415), .A2(n2416), .ZN(n15640) );
OR2_X1 U27220 ( .A1(n16450), .A2(n11362), .ZN(n2415) );
NAND2_X1 U27221 ( .A1(n16451), .A2(n2308), .ZN(n2416) );
NAND2_X1 U27222 ( .A1(n2418), .A2(n2419), .ZN(n15636) );
OR2_X1 U27223 ( .A1(n16450), .A2(n11358), .ZN(n2418) );
NAND2_X1 U27224 ( .A1(n16451), .A2(n2051), .ZN(n2419) );
NAND2_X1 U27225 ( .A1(n2420), .A2(n2421), .ZN(n15634) );
OR2_X1 U27226 ( .A1(n16451), .A2(n11356), .ZN(n2420) );
NAND2_X1 U27227 ( .A1(n16452), .A2(n2018), .ZN(n2421) );
NAND2_X1 U27228 ( .A1(n2422), .A2(n2423), .ZN(n15632) );
OR2_X1 U27229 ( .A1(n16452), .A2(n11354), .ZN(n2422) );
NAND2_X1 U27230 ( .A1(n16453), .A2(n2136), .ZN(n2423) );
NAND2_X1 U27231 ( .A1(n2424), .A2(n2425), .ZN(n15630) );
OR2_X1 U27232 ( .A1(n16453), .A2(n11352), .ZN(n2424) );
NAND2_X1 U27233 ( .A1(n16450), .A2(n2426), .ZN(n2425) );
NAND2_X1 U27234 ( .A1(n2428), .A2(n2429), .ZN(n15626) );
OR2_X1 U27235 ( .A1(n16453), .A2(n11348), .ZN(n2428) );
NAND2_X1 U27236 ( .A1(n16451), .A2(n2043), .ZN(n2429) );
NAND2_X1 U27237 ( .A1(n2430), .A2(n2431), .ZN(n15624) );
OR2_X1 U27238 ( .A1(n16450), .A2(n11346), .ZN(n2430) );
NAND2_X1 U27239 ( .A1(n16451), .A2(n2432), .ZN(n2431) );
NAND2_X1 U27240 ( .A1(n1993), .A2(n1994), .ZN(n15568) );
OR2_X1 U27241 ( .A1(n16451), .A2(n11307), .ZN(n1993) );
NAND2_X1 U27242 ( .A1(n16451), .A2(crash_dump_o_75_), .ZN(n1994) );
NAND2_X1 U27243 ( .A1(n2000), .A2(n2001), .ZN(n15562) );
OR2_X1 U27244 ( .A1(n2003), .A2(n11519), .ZN(n2000) );
NAND2_X1 U27245 ( .A1(n16451), .A2(n16439), .ZN(n2001) );
NAND2_X1 U27246 ( .A1(n7287), .A2(n7288), .ZN(n15571) );
OR2_X1 U27247 ( .A1(n19973), .A2(n11309), .ZN(n7288) );
NAND2_X1 U27248 ( .A1(n19973), .A2(n7185), .ZN(n7287) );
NAND2_X1 U27249 ( .A1(n1913), .A2(n1914), .ZN(n15774) );
OR2_X1 U27250 ( .A1(n1885), .A2(n11505), .ZN(n1913) );
NAND2_X1 U27251 ( .A1(n16453), .A2(crash_dump_o_94_), .ZN(n1914) );
NAND2_X1 U27252 ( .A1(n1951), .A2(n1952), .ZN(n15769) );
OR2_X1 U27253 ( .A1(n16451), .A2(n11495), .ZN(n1951) );
NAND2_X1 U27254 ( .A1(n16453), .A2(crash_dump_o_85_), .ZN(n1952) );
NAND2_X1 U27255 ( .A1(n1910), .A2(n1911), .ZN(n15746) );
OR2_X1 U27256 ( .A1(n16452), .A2(n11467), .ZN(n1910) );
NAND2_X1 U27257 ( .A1(n16453), .A2(crash_dump_o_95_), .ZN(n1911) );
NAND2_X1 U27258 ( .A1(n1901), .A2(n1902), .ZN(n15745) );
OR2_X1 U27259 ( .A1(n1885), .A2(n11466), .ZN(n1901) );
NAND2_X1 U27260 ( .A1(n16453), .A2(crash_dump_o_69_), .ZN(n1902) );
NAND2_X1 U27261 ( .A1(n1904), .A2(n1905), .ZN(n14948) );
OR2_X1 U27262 ( .A1(n1885), .A2(n10704), .ZN(n1904) );
NAND2_X1 U27263 ( .A1(n16453), .A2(crash_dump_o_68_), .ZN(n1905) );
NAND2_X1 U27264 ( .A1(n1907), .A2(n1908), .ZN(n14914) );
OR2_X1 U27265 ( .A1(n1885), .A2(n10670), .ZN(n1907) );
NAND2_X1 U27266 ( .A1(n16453), .A2(crash_dump_o_67_), .ZN(n1908) );
NAND2_X1 U27267 ( .A1(n1916), .A2(n1917), .ZN(n14906) );
OR2_X1 U27268 ( .A1(n16450), .A2(n10662), .ZN(n1916) );
NAND2_X1 U27269 ( .A1(n16453), .A2(crash_dump_o_66_), .ZN(n1917) );
NAND2_X1 U27270 ( .A1(n2741), .A2(n2742), .ZN(n15654) );
OR2_X1 U27271 ( .A1(n1885), .A2(n11520), .ZN(n2741) );
NAND2_X1 U27272 ( .A1(n16452), .A2(n2743), .ZN(n2742) );
NAND2_X1 U27273 ( .A1(n2744), .A2(n2745), .ZN(n2743) );
AND2_X1 U27274 ( .A1(n3556), .A2(n19885), .ZN(n3061) );
NOR2_X1 U27275 ( .A1(n11459), .A2(n15812), .ZN(n3556) );
NAND2_X1 U27276 ( .A1(n5423), .A2(n5424), .ZN(n15534) );
NAND2_X1 U27277 ( .A1(n16415), .A2(n16154), .ZN(n5424) );
NOR2_X1 U27278 ( .A1(n5426), .A2(n5427), .ZN(n5423) );
NAND2_X1 U27279 ( .A1(n5428), .A2(n5429), .ZN(n15533) );
NAND2_X1 U27280 ( .A1(n5382), .A2(n16155), .ZN(n5429) );
NOR2_X1 U27281 ( .A1(n5431), .A2(n5432), .ZN(n5428) );
NAND2_X1 U27282 ( .A1(n5433), .A2(n5434), .ZN(n15532) );
NAND2_X1 U27283 ( .A1(n16415), .A2(n16156), .ZN(n5434) );
NOR2_X1 U27284 ( .A1(n5436), .A2(n5437), .ZN(n5433) );
NAND2_X1 U27285 ( .A1(n5446), .A2(n5447), .ZN(n15529) );
NAND2_X1 U27286 ( .A1(n5382), .A2(n16157), .ZN(n5447) );
NOR2_X1 U27287 ( .A1(n5449), .A2(n5450), .ZN(n5446) );
NAND2_X1 U27288 ( .A1(n5475), .A2(n5476), .ZN(n15522) );
NAND2_X1 U27289 ( .A1(n5382), .A2(n16158), .ZN(n5476) );
NOR2_X1 U27290 ( .A1(n5478), .A2(n5479), .ZN(n5475) );
NAND2_X1 U27291 ( .A1(n5480), .A2(n5481), .ZN(n15521) );
NAND2_X1 U27292 ( .A1(n5382), .A2(n16159), .ZN(n5481) );
NOR2_X1 U27293 ( .A1(n5483), .A2(n5484), .ZN(n5480) );
NAND2_X1 U27294 ( .A1(n5485), .A2(n5486), .ZN(n15520) );
NAND2_X1 U27295 ( .A1(n5382), .A2(n16160), .ZN(n5486) );
NOR2_X1 U27296 ( .A1(n5488), .A2(n5489), .ZN(n5485) );
NAND2_X1 U27297 ( .A1(n5490), .A2(n5491), .ZN(n15519) );
NAND2_X1 U27298 ( .A1(n5382), .A2(n16161), .ZN(n5491) );
NOR2_X1 U27299 ( .A1(n5493), .A2(n5494), .ZN(n5490) );
NAND2_X1 U27300 ( .A1(n5495), .A2(n5496), .ZN(n15518) );
NAND2_X1 U27301 ( .A1(n16415), .A2(n16162), .ZN(n5496) );
NOR2_X1 U27302 ( .A1(n5498), .A2(n5499), .ZN(n5495) );
NAND2_X1 U27303 ( .A1(n5500), .A2(n5501), .ZN(n15517) );
NAND2_X1 U27304 ( .A1(n5382), .A2(n16163), .ZN(n5501) );
NOR2_X1 U27305 ( .A1(n5503), .A2(n5504), .ZN(n5500) );
NAND2_X1 U27306 ( .A1(n5513), .A2(n5514), .ZN(n15514) );
NAND2_X1 U27307 ( .A1(n16415), .A2(n16164), .ZN(n5514) );
NOR2_X1 U27308 ( .A1(n5516), .A2(n5517), .ZN(n5513) );
NAND2_X1 U27309 ( .A1(n5518), .A2(n5519), .ZN(n15513) );
NAND2_X1 U27310 ( .A1(n5382), .A2(n16165), .ZN(n5519) );
NOR2_X1 U27311 ( .A1(n5521), .A2(n5522), .ZN(n5518) );
NAND2_X1 U27312 ( .A1(n5523), .A2(n5524), .ZN(n15512) );
NAND2_X1 U27313 ( .A1(n16415), .A2(n16166), .ZN(n5524) );
NOR2_X1 U27314 ( .A1(n5526), .A2(n5527), .ZN(n5523) );
NAND2_X1 U27315 ( .A1(n4116), .A2(n4117), .ZN(n15496) );
NAND2_X1 U27316 ( .A1(n4061), .A2(n16167), .ZN(n4117) );
NOR2_X1 U27317 ( .A1(n4119), .A2(n4120), .ZN(n4116) );
NAND2_X1 U27318 ( .A1(n4182), .A2(n4183), .ZN(n15485) );
NAND2_X1 U27319 ( .A1(n16427), .A2(n16168), .ZN(n4183) );
NOR2_X1 U27320 ( .A1(n4185), .A2(n4186), .ZN(n4182) );
NAND2_X1 U27321 ( .A1(n4236), .A2(n4237), .ZN(n15476) );
NAND2_X1 U27322 ( .A1(n16427), .A2(n16169), .ZN(n4237) );
NOR2_X1 U27323 ( .A1(n4239), .A2(n4240), .ZN(n4236) );
NAND2_X1 U27324 ( .A1(n4242), .A2(n4243), .ZN(n15475) );
NAND2_X1 U27325 ( .A1(n16427), .A2(n16170), .ZN(n4243) );
NOR2_X1 U27326 ( .A1(n4245), .A2(n4246), .ZN(n4242) );
NAND2_X1 U27327 ( .A1(n4248), .A2(n4249), .ZN(n15474) );
NAND2_X1 U27328 ( .A1(n16427), .A2(n16171), .ZN(n4249) );
NOR2_X1 U27329 ( .A1(n4253), .A2(n4254), .ZN(n4248) );
NAND2_X1 U27330 ( .A1(n5301), .A2(n5302), .ZN(n15462) );
NAND2_X1 U27331 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_30), .ZN(n5302) );
NAND2_X1 U27332 ( .A1(n5278), .A2(n16172), .ZN(n5301) );
NAND2_X1 U27333 ( .A1(n5304), .A2(n5305), .ZN(n15461) );
NAND2_X1 U27334 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_2), .ZN(n5305) );
NAND2_X1 U27335 ( .A1(n5278), .A2(n16173), .ZN(n5304) );
NAND2_X1 U27336 ( .A1(n5307), .A2(n5308), .ZN(n15460) );
NAND2_X1 U27337 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_29), .ZN(n5308) );
NAND2_X1 U27338 ( .A1(n16416), .A2(n16174), .ZN(n5307) );
NAND2_X1 U27339 ( .A1(n5310), .A2(n5311), .ZN(n15459) );
NAND2_X1 U27340 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_28), .ZN(n5311) );
NAND2_X1 U27341 ( .A1(n5278), .A2(n16175), .ZN(n5310) );
NAND2_X1 U27342 ( .A1(n5313), .A2(n5314), .ZN(n15458) );
NAND2_X1 U27343 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_27), .ZN(n5314) );
NAND2_X1 U27344 ( .A1(n16416), .A2(n16176), .ZN(n5313) );
NAND2_X1 U27345 ( .A1(n5316), .A2(n5317), .ZN(n15457) );
NAND2_X1 U27346 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_26), .ZN(n5317) );
NAND2_X1 U27347 ( .A1(n5278), .A2(n16177), .ZN(n5316) );
NAND2_X1 U27348 ( .A1(n5319), .A2(n5320), .ZN(n15456) );
NAND2_X1 U27349 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_25), .ZN(n5320) );
NAND2_X1 U27350 ( .A1(n16416), .A2(n16178), .ZN(n5319) );
NAND2_X1 U27351 ( .A1(n5322), .A2(n5323), .ZN(n15455) );
NAND2_X1 U27352 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_24), .ZN(n5323) );
NAND2_X1 U27353 ( .A1(n5278), .A2(n16179), .ZN(n5322) );
NAND2_X1 U27354 ( .A1(n5325), .A2(n5326), .ZN(n15454) );
NAND2_X1 U27355 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_23), .ZN(n5326) );
NAND2_X1 U27356 ( .A1(n16416), .A2(n16180), .ZN(n5325) );
NAND2_X1 U27357 ( .A1(n5328), .A2(n5329), .ZN(n15453) );
NAND2_X1 U27358 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_22), .ZN(n5329) );
NAND2_X1 U27359 ( .A1(n5278), .A2(n16181), .ZN(n5328) );
NAND2_X1 U27360 ( .A1(n5331), .A2(n5332), .ZN(n15452) );
NAND2_X1 U27361 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_21), .ZN(n5332) );
NAND2_X1 U27362 ( .A1(n16416), .A2(n16182), .ZN(n5331) );
NAND2_X1 U27363 ( .A1(n5334), .A2(n5335), .ZN(n15451) );
NAND2_X1 U27364 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_20), .ZN(n5335) );
NAND2_X1 U27365 ( .A1(n5278), .A2(n16183), .ZN(n5334) );
NAND2_X1 U27366 ( .A1(n5337), .A2(n5338), .ZN(n15450) );
NAND2_X1 U27367 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_1), .ZN(n5338) );
NAND2_X1 U27368 ( .A1(n5278), .A2(n16184), .ZN(n5337) );
NAND2_X1 U27369 ( .A1(n5340), .A2(n5341), .ZN(n15449) );
NAND2_X1 U27370 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_19), .ZN(n5341) );
NAND2_X1 U27371 ( .A1(n5278), .A2(n16185), .ZN(n5340) );
NAND2_X1 U27372 ( .A1(n5343), .A2(n5344), .ZN(n15448) );
NAND2_X1 U27373 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_18), .ZN(n5344) );
NAND2_X1 U27374 ( .A1(n5278), .A2(n16186), .ZN(n5343) );
NAND2_X1 U27375 ( .A1(n5346), .A2(n5347), .ZN(n15447) );
NAND2_X1 U27376 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_17), .ZN(n5347) );
NAND2_X1 U27377 ( .A1(n5278), .A2(n16187), .ZN(n5346) );
NAND2_X1 U27378 ( .A1(n5349), .A2(n5350), .ZN(n15446) );
NAND2_X1 U27379 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_16), .ZN(n5350) );
NAND2_X1 U27380 ( .A1(n5278), .A2(n16188), .ZN(n5349) );
NAND2_X1 U27381 ( .A1(n5352), .A2(n5353), .ZN(n15445) );
NAND2_X1 U27382 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_15), .ZN(n5353) );
NAND2_X1 U27383 ( .A1(n5278), .A2(n16189), .ZN(n5352) );
NAND2_X1 U27384 ( .A1(n5355), .A2(n5356), .ZN(n15444) );
NAND2_X1 U27385 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_14), .ZN(n5356) );
NAND2_X1 U27386 ( .A1(n16416), .A2(n16190), .ZN(n5355) );
NAND2_X1 U27387 ( .A1(n5358), .A2(n5359), .ZN(n15443) );
NAND2_X1 U27388 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_13), .ZN(n5359) );
NAND2_X1 U27389 ( .A1(n5278), .A2(n16191), .ZN(n5358) );
NAND2_X1 U27390 ( .A1(n5361), .A2(n5362), .ZN(n15442) );
NAND2_X1 U27391 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_12), .ZN(n5362) );
NAND2_X1 U27392 ( .A1(n16416), .A2(n16192), .ZN(n5361) );
NAND2_X1 U27393 ( .A1(n5364), .A2(n5365), .ZN(n15421) );
NAND2_X1 U27394 ( .A1(n5277), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_11), .ZN(n5365) );
NAND2_X1 U27395 ( .A1(n5278), .A2(n16193), .ZN(n5364) );
NAND2_X1 U27396 ( .A1(n5367), .A2(n5368), .ZN(n15420) );
NAND2_X1 U27397 ( .A1(n16417), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_one_shift_10), .ZN(n5368) );
NAND2_X1 U27398 ( .A1(n16416), .A2(n16194), .ZN(n5367) );
NAND2_X1 U27399 ( .A1(n7807), .A2(n7808), .ZN(n15363) );
OR2_X1 U27400 ( .A1(n19977), .A2(n11110), .ZN(n7807) );
NAND2_X1 U27401 ( .A1(n16348), .A2(n7191), .ZN(n7808) );
NAND2_X1 U27402 ( .A1(n7805), .A2(n7806), .ZN(n14958) );
OR2_X1 U27403 ( .A1(n16349), .A2(n10714), .ZN(n7805) );
NAND2_X1 U27404 ( .A1(n16348), .A2(n7188), .ZN(n7806) );
NAND2_X1 U27405 ( .A1(n2990), .A2(n2991), .ZN(n14822) );
NAND2_X1 U27406 ( .A1(n2897), .A2(n16052), .ZN(n2991) );
NOR2_X1 U27407 ( .A1(n2992), .A2(n2993), .ZN(n2990) );
NOR2_X1 U27408 ( .A1(n10580), .A2(n16444), .ZN(n2992) );
NAND2_X1 U27409 ( .A1(n2974), .A2(n2975), .ZN(n14814) );
NAND2_X1 U27410 ( .A1(n16445), .A2(n16053), .ZN(n2975) );
NOR2_X1 U27411 ( .A1(n2976), .A2(n2977), .ZN(n2974) );
NOR2_X1 U27412 ( .A1(n10572), .A2(n2900), .ZN(n2976) );
NAND2_X1 U27413 ( .A1(n2954), .A2(n2955), .ZN(n14804) );
NAND2_X1 U27414 ( .A1(n2897), .A2(n16054), .ZN(n2955) );
NOR2_X1 U27415 ( .A1(n2956), .A2(n2957), .ZN(n2954) );
NOR2_X1 U27416 ( .A1(n10562), .A2(n16444), .ZN(n2956) );
NAND2_X1 U27417 ( .A1(n2946), .A2(n2947), .ZN(n14800) );
NAND2_X1 U27418 ( .A1(n16445), .A2(n16055), .ZN(n2947) );
NOR2_X1 U27419 ( .A1(n2948), .A2(n2949), .ZN(n2946) );
NOR2_X1 U27420 ( .A1(n10558), .A2(n16444), .ZN(n2948) );
NAND2_X1 U27421 ( .A1(n2942), .A2(n2943), .ZN(n14798) );
NAND2_X1 U27422 ( .A1(n2897), .A2(n16056), .ZN(n2943) );
NOR2_X1 U27423 ( .A1(n2944), .A2(n2945), .ZN(n2942) );
NOR2_X1 U27424 ( .A1(n10556), .A2(n2900), .ZN(n2944) );
NAND2_X1 U27425 ( .A1(n1634), .A2(n1635), .ZN(n15309) );
OR2_X1 U27426 ( .A1(n16460), .A2(n11492), .ZN(n1635) );
NAND2_X1 U27427 ( .A1(data_addr_o_29_), .A2(n16460), .ZN(n1634) );
NAND2_X1 U27428 ( .A1(n1636), .A2(n1637), .ZN(n15308) );
OR2_X1 U27429 ( .A1(n16460), .A2(n11058), .ZN(n1637) );
NAND2_X1 U27430 ( .A1(data_addr_o_28_), .A2(n1606), .ZN(n1636) );
NAND2_X1 U27431 ( .A1(n1638), .A2(n1639), .ZN(n15307) );
OR2_X1 U27432 ( .A1(n16460), .A2(n11057), .ZN(n1639) );
NAND2_X1 U27433 ( .A1(data_addr_o_27_), .A2(n16460), .ZN(n1638) );
NAND2_X1 U27434 ( .A1(n1640), .A2(n1641), .ZN(n15306) );
OR2_X1 U27435 ( .A1(n16460), .A2(n11056), .ZN(n1641) );
NAND2_X1 U27436 ( .A1(data_addr_o_26_), .A2(n16460), .ZN(n1640) );
NAND2_X1 U27437 ( .A1(n1642), .A2(n1643), .ZN(n15305) );
OR2_X1 U27438 ( .A1(n16460), .A2(n11055), .ZN(n1643) );
NAND2_X1 U27439 ( .A1(data_addr_o_25_), .A2(n16460), .ZN(n1642) );
NAND2_X1 U27440 ( .A1(n1644), .A2(n1645), .ZN(n15304) );
OR2_X1 U27441 ( .A1(n16460), .A2(n11054), .ZN(n1645) );
NAND2_X1 U27442 ( .A1(data_addr_o_24_), .A2(n1606), .ZN(n1644) );
NAND2_X1 U27443 ( .A1(n1646), .A2(n1647), .ZN(n15303) );
OR2_X1 U27444 ( .A1(n16460), .A2(n11053), .ZN(n1647) );
NAND2_X1 U27445 ( .A1(data_addr_o_23_), .A2(n1606), .ZN(n1646) );
NAND2_X1 U27446 ( .A1(n1648), .A2(n1649), .ZN(n15302) );
OR2_X1 U27447 ( .A1(n16460), .A2(n11052), .ZN(n1649) );
NAND2_X1 U27448 ( .A1(data_addr_o_22_), .A2(n16460), .ZN(n1648) );
NAND2_X1 U27449 ( .A1(n1653), .A2(n1654), .ZN(n15300) );
OR2_X1 U27450 ( .A1(n16460), .A2(n11050), .ZN(n1654) );
NAND2_X1 U27451 ( .A1(data_addr_o_20_), .A2(n1606), .ZN(n1653) );
NAND2_X1 U27452 ( .A1(n1659), .A2(n1660), .ZN(n15299) );
OR2_X1 U27453 ( .A1(n16460), .A2(n11049), .ZN(n1660) );
NAND2_X1 U27454 ( .A1(data_addr_o_19_), .A2(n1606), .ZN(n1659) );
NAND2_X1 U27455 ( .A1(n1661), .A2(n1662), .ZN(n15298) );
OR2_X1 U27456 ( .A1(n16460), .A2(n11048), .ZN(n1662) );
NAND2_X1 U27457 ( .A1(data_addr_o_18_), .A2(n1606), .ZN(n1661) );
NAND2_X1 U27458 ( .A1(n1663), .A2(n1664), .ZN(n15297) );
OR2_X1 U27459 ( .A1(n16460), .A2(n11047), .ZN(n1664) );
NAND2_X1 U27460 ( .A1(data_addr_o_17_), .A2(n1606), .ZN(n1663) );
NAND2_X1 U27461 ( .A1(n1665), .A2(n1666), .ZN(n15296) );
OR2_X1 U27462 ( .A1(n16460), .A2(n11046), .ZN(n1666) );
NAND2_X1 U27463 ( .A1(data_addr_o_16_), .A2(n1606), .ZN(n1665) );
NAND2_X1 U27464 ( .A1(n5662), .A2(n5663), .ZN(n15510) );
NAND2_X1 U27465 ( .A1(n11256), .A2(n20906), .ZN(n5663) );
NOR2_X1 U27466 ( .A1(n5651), .A2(n5664), .ZN(n5662) );
NOR2_X1 U27467 ( .A1(n11256), .A2(n20906), .ZN(n5664) );
NAND2_X1 U27468 ( .A1(n5659), .A2(n5660), .ZN(n15509) );
NAND2_X1 U27469 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N218), .A2(n20906), .ZN(n5660) );
NOR2_X1 U27470 ( .A1(n5651), .A2(n5661), .ZN(n5659) );
NOR2_X1 U27471 ( .A1(n11255), .A2(n20906), .ZN(n5661) );
NAND2_X1 U27472 ( .A1(n5656), .A2(n5657), .ZN(n15508) );
NAND2_X1 U27473 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N219), .A2(n20906), .ZN(n5657) );
NOR2_X1 U27474 ( .A1(n5651), .A2(n5658), .ZN(n5656) );
NOR2_X1 U27475 ( .A1(n11254), .A2(n20906), .ZN(n5658) );
NAND2_X1 U27476 ( .A1(n5653), .A2(n5654), .ZN(n15507) );
NAND2_X1 U27477 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N220), .A2(n20906), .ZN(n5654) );
NOR2_X1 U27478 ( .A1(n5651), .A2(n5655), .ZN(n5653) );
NOR2_X1 U27479 ( .A1(n11253), .A2(n20906), .ZN(n5655) );
NAND2_X1 U27480 ( .A1(n5649), .A2(n5650), .ZN(n15506) );
NAND2_X1 U27481 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_N221), .A2(n20906), .ZN(n5650) );
NOR2_X1 U27482 ( .A1(n5651), .A2(n5652), .ZN(n5649) );
NOR2_X1 U27483 ( .A1(n11252), .A2(n20906), .ZN(n5652) );
INV_X1 U27484 ( .A(rst_ni), .ZN(n19748) );
NAND2_X1 U27485 ( .A1(n4413), .A2(n4414), .ZN(n15408) );
NAND2_X1 U27486 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_32), .A2(n20909), .ZN(n4414) );
NOR2_X1 U27487 ( .A1(n4415), .A2(n4416), .ZN(n4413) );
NOR2_X1 U27488 ( .A1(n11154), .A2(n4410), .ZN(n4416) );
NAND2_X1 U27489 ( .A1(n4406), .A2(n4407), .ZN(n15407) );
NAND2_X1 U27490 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_33), .A2(n20909), .ZN(n4407) );
NOR2_X1 U27491 ( .A1(n4408), .A2(n4409), .ZN(n4406) );
NOR2_X1 U27492 ( .A1(n11153), .A2(n4410), .ZN(n4409) );
NAND2_X1 U27493 ( .A1(n8084), .A2(n8085), .ZN(n15025) );
NAND2_X1 U27494 ( .A1(n20988), .A2(priv_mode_id_1), .ZN(n8085) );
NOR2_X1 U27495 ( .A1(n8086), .A2(n8087), .ZN(n8084) );
NOR2_X1 U27496 ( .A1(n10780), .A2(n8074), .ZN(n8087) );
NAND2_X1 U27497 ( .A1(n8123), .A2(n8124), .ZN(n15021) );
NAND2_X1 U27498 ( .A1(n20988), .A2(priv_mode_id_0), .ZN(n8124) );
NOR2_X1 U27499 ( .A1(n8086), .A2(n8125), .ZN(n8123) );
NOR2_X1 U27500 ( .A1(n11303), .A2(n8074), .ZN(n8125) );
NAND2_X1 U27501 ( .A1(n8075), .A2(n8076), .ZN(n15020) );
OR2_X1 U27502 ( .A1(n20988), .A2(n10777), .ZN(n8075) );
NAND2_X1 U27503 ( .A1(n20988), .A2(n8077), .ZN(n8076) );
NAND2_X1 U27504 ( .A1(n15909), .A2(n8078), .ZN(n8077) );
NAND2_X1 U27505 ( .A1(n5666), .A2(n5667), .ZN(n15473) );
OR2_X1 U27506 ( .A1(n5668), .A2(n11219), .ZN(n5666) );
NAND2_X1 U27507 ( .A1(n5668), .A2(ex_block_i_alu_is_equal_result), .ZN(n5667) );
NOR2_X1 U27508 ( .A1(n4411), .A2(n5374), .ZN(n5668) );
NAND2_X1 U27509 ( .A1(n3034), .A2(n3035), .ZN(n15740) );
NAND2_X1 U27510 ( .A1(n19885), .A2(n3036), .ZN(n3035) );
NOR2_X1 U27511 ( .A1(n3037), .A2(n3038), .ZN(n3034) );
NOR2_X1 U27512 ( .A1(n11459), .A2(n3039), .ZN(n3038) );
NAND2_X1 U27513 ( .A1(n7224), .A2(n7225), .ZN(n15396) );
OR2_X1 U27514 ( .A1(n7178), .A2(n11143), .ZN(n7225) );
NAND2_X1 U27515 ( .A1(n7178), .A2(n7226), .ZN(n7224) );
NAND2_X1 U27516 ( .A1(n7201), .A2(n7202), .ZN(n15395) );
OR2_X1 U27517 ( .A1(n7178), .A2(n11142), .ZN(n7202) );
NAND2_X1 U27518 ( .A1(n7178), .A2(n7203), .ZN(n7201) );
NAND2_X1 U27519 ( .A1(n7246), .A2(n7247), .ZN(n15392) );
OR2_X1 U27520 ( .A1(n16398), .A2(n11139), .ZN(n7247) );
NAND2_X1 U27521 ( .A1(n16398), .A2(n7069), .ZN(n7246) );
NAND2_X1 U27522 ( .A1(n7244), .A2(n7245), .ZN(n15391) );
OR2_X1 U27523 ( .A1(n16398), .A2(n11138), .ZN(n7245) );
NAND2_X1 U27524 ( .A1(n16397), .A2(n7068), .ZN(n7244) );
NAND2_X1 U27525 ( .A1(n7220), .A2(n7221), .ZN(n15390) );
OR2_X1 U27526 ( .A1(n7178), .A2(n11137), .ZN(n7221) );
NAND2_X1 U27527 ( .A1(n16398), .A2(n6896), .ZN(n7220) );
NAND2_X1 U27528 ( .A1(n7204), .A2(n7205), .ZN(n15389) );
OR2_X1 U27529 ( .A1(n16397), .A2(n11136), .ZN(n7205) );
NAND2_X1 U27530 ( .A1(n7178), .A2(n6824), .ZN(n7204) );
NAND2_X1 U27531 ( .A1(n7197), .A2(n7198), .ZN(n15387) );
OR2_X1 U27532 ( .A1(n16398), .A2(n11134), .ZN(n7198) );
NAND2_X1 U27533 ( .A1(n7178), .A2(n6792), .ZN(n7197) );
NAND2_X1 U27534 ( .A1(n7251), .A2(n7252), .ZN(n15386) );
OR2_X1 U27535 ( .A1(n16398), .A2(n11133), .ZN(n7252) );
NAND2_X1 U27536 ( .A1(n16398), .A2(n7253), .ZN(n7251) );
NAND2_X1 U27537 ( .A1(n7840), .A2(n7841), .ZN(n15366) );
OR2_X1 U27538 ( .A1(n16349), .A2(n11113), .ZN(n7841) );
NAND2_X1 U27539 ( .A1(n16349), .A2(n7226), .ZN(n7840) );
NAND2_X1 U27540 ( .A1(n7817), .A2(n7818), .ZN(n15365) );
OR2_X1 U27541 ( .A1(n16348), .A2(n11112), .ZN(n7818) );
NAND2_X1 U27542 ( .A1(n16348), .A2(n7203), .ZN(n7817) );
NAND2_X1 U27543 ( .A1(n7811), .A2(n7812), .ZN(n15364) );
OR2_X1 U27544 ( .A1(n19977), .A2(n11111), .ZN(n7812) );
NAND2_X1 U27545 ( .A1(n16348), .A2(n7037), .ZN(n7811) );
NAND2_X1 U27546 ( .A1(n7819), .A2(n7820), .ZN(n15359) );
OR2_X1 U27547 ( .A1(n16349), .A2(n11106), .ZN(n7820) );
NAND2_X1 U27548 ( .A1(n16348), .A2(n6824), .ZN(n7819) );
NAND2_X1 U27549 ( .A1(n7815), .A2(n7816), .ZN(n15358) );
OR2_X1 U27550 ( .A1(n16348), .A2(n11105), .ZN(n7816) );
NAND2_X1 U27551 ( .A1(n16348), .A2(n6803), .ZN(n7815) );
NAND2_X1 U27552 ( .A1(n7813), .A2(n7814), .ZN(n15357) );
OR2_X1 U27553 ( .A1(n19977), .A2(n11104), .ZN(n7814) );
NAND2_X1 U27554 ( .A1(n16349), .A2(n6792), .ZN(n7813) );
NAND2_X1 U27555 ( .A1(n7864), .A2(n7865), .ZN(n15356) );
OR2_X1 U27556 ( .A1(n19977), .A2(n11103), .ZN(n7865) );
NAND2_X1 U27557 ( .A1(n16348), .A2(n7253), .ZN(n7864) );
NAND2_X1 U27558 ( .A1(n7208), .A2(n7209), .ZN(n15220) );
OR2_X1 U27559 ( .A1(n7178), .A2(n10975), .ZN(n7209) );
NAND2_X1 U27560 ( .A1(n7178), .A2(n6842), .ZN(n7208) );
NAND2_X1 U27561 ( .A1(n7823), .A2(n7824), .ZN(n15219) );
OR2_X1 U27562 ( .A1(n16349), .A2(n10974), .ZN(n7824) );
NAND2_X1 U27563 ( .A1(n16349), .A2(n6842), .ZN(n7823) );
NAND2_X1 U27564 ( .A1(n7210), .A2(n7211), .ZN(n15205) );
OR2_X1 U27565 ( .A1(n16397), .A2(n10960), .ZN(n7211) );
NAND2_X1 U27566 ( .A1(n16397), .A2(n6851), .ZN(n7210) );
NAND2_X1 U27567 ( .A1(n7825), .A2(n7826), .ZN(n15204) );
OR2_X1 U27568 ( .A1(n16348), .A2(n10959), .ZN(n7826) );
NAND2_X1 U27569 ( .A1(n16349), .A2(n6851), .ZN(n7825) );
NAND2_X1 U27570 ( .A1(n7212), .A2(n7213), .ZN(n15190) );
OR2_X1 U27571 ( .A1(n16397), .A2(n10945), .ZN(n7213) );
NAND2_X1 U27572 ( .A1(n16398), .A2(n6860), .ZN(n7212) );
NAND2_X1 U27573 ( .A1(n7827), .A2(n7828), .ZN(n15189) );
OR2_X1 U27574 ( .A1(n19977), .A2(n10944), .ZN(n7828) );
NAND2_X1 U27575 ( .A1(n16349), .A2(n6860), .ZN(n7827) );
NAND2_X1 U27576 ( .A1(n7214), .A2(n7215), .ZN(n15175) );
OR2_X1 U27577 ( .A1(n16398), .A2(n10930), .ZN(n7215) );
NAND2_X1 U27578 ( .A1(n16398), .A2(n6869), .ZN(n7214) );
NAND2_X1 U27579 ( .A1(n7829), .A2(n7830), .ZN(n15174) );
OR2_X1 U27580 ( .A1(n16348), .A2(n10929), .ZN(n7830) );
NAND2_X1 U27581 ( .A1(n16349), .A2(n6869), .ZN(n7829) );
NAND2_X1 U27582 ( .A1(n7216), .A2(n7217), .ZN(n15160) );
OR2_X1 U27583 ( .A1(n16397), .A2(n10915), .ZN(n7217) );
NAND2_X1 U27584 ( .A1(n7178), .A2(n6878), .ZN(n7216) );
NAND2_X1 U27585 ( .A1(n7831), .A2(n7832), .ZN(n15159) );
OR2_X1 U27586 ( .A1(n19977), .A2(n10914), .ZN(n7832) );
NAND2_X1 U27587 ( .A1(n16349), .A2(n6878), .ZN(n7831) );
NAND2_X1 U27588 ( .A1(n7218), .A2(n7219), .ZN(n15145) );
OR2_X1 U27589 ( .A1(n7178), .A2(n10900), .ZN(n7219) );
NAND2_X1 U27590 ( .A1(n16397), .A2(n6887), .ZN(n7218) );
NAND2_X1 U27591 ( .A1(n7833), .A2(n7834), .ZN(n15144) );
OR2_X1 U27592 ( .A1(n16349), .A2(n10899), .ZN(n7834) );
NAND2_X1 U27593 ( .A1(n16349), .A2(n6887), .ZN(n7833) );
NAND2_X1 U27594 ( .A1(n7222), .A2(n7223), .ZN(n15130) );
OR2_X1 U27595 ( .A1(n16398), .A2(n10885), .ZN(n7223) );
NAND2_X1 U27596 ( .A1(n7178), .A2(n6905), .ZN(n7222) );
NAND2_X1 U27597 ( .A1(n7838), .A2(n7839), .ZN(n15129) );
OR2_X1 U27598 ( .A1(n16349), .A2(n10884), .ZN(n7839) );
NAND2_X1 U27599 ( .A1(n16349), .A2(n6905), .ZN(n7838) );
NAND2_X1 U27600 ( .A1(n7227), .A2(n7228), .ZN(n15115) );
OR2_X1 U27601 ( .A1(n7178), .A2(n10870), .ZN(n7228) );
NAND2_X1 U27602 ( .A1(n16398), .A2(n6925), .ZN(n7227) );
NAND2_X1 U27603 ( .A1(n7229), .A2(n7230), .ZN(n15098) );
OR2_X1 U27604 ( .A1(n16398), .A2(n10853), .ZN(n7230) );
NAND2_X1 U27605 ( .A1(n16397), .A2(n6934), .ZN(n7229) );
NAND2_X1 U27606 ( .A1(n7844), .A2(n7845), .ZN(n15097) );
OR2_X1 U27607 ( .A1(n16348), .A2(n10852), .ZN(n7845) );
NAND2_X1 U27608 ( .A1(n16349), .A2(n6934), .ZN(n7844) );
NAND2_X1 U27609 ( .A1(n7233), .A2(n7234), .ZN(n15083) );
OR2_X1 U27610 ( .A1(n7178), .A2(n10838), .ZN(n7234) );
NAND2_X1 U27611 ( .A1(n7178), .A2(n6952), .ZN(n7233) );
NAND2_X1 U27612 ( .A1(n7235), .A2(n7236), .ZN(n15069) );
OR2_X1 U27613 ( .A1(n16398), .A2(n10824), .ZN(n7236) );
NAND2_X1 U27614 ( .A1(n16398), .A2(n7237), .ZN(n7235) );
NAND2_X1 U27615 ( .A1(n7238), .A2(n7239), .ZN(n15054) );
OR2_X1 U27616 ( .A1(n7178), .A2(n10809), .ZN(n7239) );
NAND2_X1 U27617 ( .A1(n16397), .A2(n7240), .ZN(n7238) );
NAND2_X1 U27618 ( .A1(n7241), .A2(n7242), .ZN(n15040) );
OR2_X1 U27619 ( .A1(n16398), .A2(n10795), .ZN(n7242) );
NAND2_X1 U27620 ( .A1(n7178), .A2(n7243), .ZN(n7241) );
NAND2_X1 U27621 ( .A1(n7248), .A2(n7249), .ZN(n15001) );
OR2_X1 U27622 ( .A1(n16398), .A2(n10757), .ZN(n7249) );
NAND2_X1 U27623 ( .A1(n16398), .A2(n7250), .ZN(n7248) );
NAND2_X1 U27624 ( .A1(n7796), .A2(n7797), .ZN(n14986) );
OR2_X1 U27625 ( .A1(n16348), .A2(n10742), .ZN(n7797) );
NAND2_X1 U27626 ( .A1(n16348), .A2(n7179), .ZN(n7796) );
NAND2_X1 U27627 ( .A1(n7799), .A2(n7800), .ZN(n14972) );
OR2_X1 U27628 ( .A1(n19977), .A2(n10728), .ZN(n7800) );
NAND2_X1 U27629 ( .A1(n16348), .A2(n7182), .ZN(n7799) );
NAND2_X1 U27630 ( .A1(n7809), .A2(n7810), .ZN(n14945) );
OR2_X1 U27631 ( .A1(n19977), .A2(n10701), .ZN(n7810) );
NAND2_X1 U27632 ( .A1(n16348), .A2(n7194), .ZN(n7809) );
NAND2_X1 U27633 ( .A1(n7231), .A2(n7232), .ZN(n14903) );
OR2_X1 U27634 ( .A1(n16398), .A2(n10659), .ZN(n7232) );
NAND2_X1 U27635 ( .A1(n16397), .A2(n6943), .ZN(n7231) );
NAND2_X1 U27636 ( .A1(n7206), .A2(n7207), .ZN(n14885) );
OR2_X1 U27637 ( .A1(n16397), .A2(n10642), .ZN(n7207) );
NAND2_X1 U27638 ( .A1(n16397), .A2(n6833), .ZN(n7206) );
NAND2_X1 U27639 ( .A1(n7821), .A2(n7822), .ZN(n14884) );
OR2_X1 U27640 ( .A1(n16349), .A2(n10641), .ZN(n7822) );
NAND2_X1 U27641 ( .A1(n16348), .A2(n6833), .ZN(n7821) );
NAND2_X1 U27642 ( .A1(n1454), .A2(n1455), .ZN(n15340) );
NAND2_X1 U27643 ( .A1(n1452), .A2(n16057), .ZN(n1455) );
NAND2_X1 U27644 ( .A1(n16465), .A2(data_rdata_i_8_), .ZN(n1454) );
NAND2_X1 U27645 ( .A1(n1456), .A2(n1457), .ZN(n15339) );
NAND2_X1 U27646 ( .A1(n1452), .A2(n16058), .ZN(n1457) );
NAND2_X1 U27647 ( .A1(n16465), .A2(data_rdata_i_31_), .ZN(n1456) );
NAND2_X1 U27648 ( .A1(n1458), .A2(n1459), .ZN(n15338) );
NAND2_X1 U27649 ( .A1(n1452), .A2(n16059), .ZN(n1459) );
NAND2_X1 U27650 ( .A1(n16465), .A2(data_rdata_i_30_), .ZN(n1458) );
NAND2_X1 U27651 ( .A1(n1460), .A2(n1461), .ZN(n15337) );
NAND2_X1 U27652 ( .A1(n1452), .A2(n16060), .ZN(n1461) );
NAND2_X1 U27653 ( .A1(n16465), .A2(data_rdata_i_29_), .ZN(n1460) );
NAND2_X1 U27654 ( .A1(n1462), .A2(n1463), .ZN(n15336) );
NAND2_X1 U27655 ( .A1(n1452), .A2(n16061), .ZN(n1463) );
NAND2_X1 U27656 ( .A1(n16465), .A2(data_rdata_i_28_), .ZN(n1462) );
NAND2_X1 U27657 ( .A1(n1464), .A2(n1465), .ZN(n15335) );
NAND2_X1 U27658 ( .A1(n1452), .A2(n16062), .ZN(n1465) );
NAND2_X1 U27659 ( .A1(n16465), .A2(data_rdata_i_27_), .ZN(n1464) );
NAND2_X1 U27660 ( .A1(n1466), .A2(n1467), .ZN(n15334) );
NAND2_X1 U27661 ( .A1(n1452), .A2(n16063), .ZN(n1467) );
NAND2_X1 U27662 ( .A1(n16465), .A2(data_rdata_i_26_), .ZN(n1466) );
NAND2_X1 U27663 ( .A1(n1468), .A2(n1469), .ZN(n15333) );
NAND2_X1 U27664 ( .A1(n1452), .A2(n16064), .ZN(n1469) );
NAND2_X1 U27665 ( .A1(n16465), .A2(data_rdata_i_25_), .ZN(n1468) );
NAND2_X1 U27666 ( .A1(n1470), .A2(n1471), .ZN(n15332) );
NAND2_X1 U27667 ( .A1(n1452), .A2(n16065), .ZN(n1471) );
NAND2_X1 U27668 ( .A1(n16465), .A2(data_rdata_i_24_), .ZN(n1470) );
NAND2_X1 U27669 ( .A1(n1472), .A2(n1473), .ZN(n15331) );
NAND2_X1 U27670 ( .A1(n1452), .A2(n16066), .ZN(n1473) );
NAND2_X1 U27671 ( .A1(n16465), .A2(data_rdata_i_23_), .ZN(n1472) );
NAND2_X1 U27672 ( .A1(n1474), .A2(n1475), .ZN(n15330) );
NAND2_X1 U27673 ( .A1(n1452), .A2(n16067), .ZN(n1475) );
NAND2_X1 U27674 ( .A1(n16465), .A2(data_rdata_i_22_), .ZN(n1474) );
NAND2_X1 U27675 ( .A1(n1476), .A2(n1477), .ZN(n15329) );
NAND2_X1 U27676 ( .A1(n1452), .A2(n16068), .ZN(n1477) );
NAND2_X1 U27677 ( .A1(n16465), .A2(data_rdata_i_21_), .ZN(n1476) );
NAND2_X1 U27678 ( .A1(n1478), .A2(n1479), .ZN(n15328) );
NAND2_X1 U27679 ( .A1(n1452), .A2(n16069), .ZN(n1479) );
NAND2_X1 U27680 ( .A1(n16465), .A2(data_rdata_i_20_), .ZN(n1478) );
NAND2_X1 U27681 ( .A1(n1480), .A2(n1481), .ZN(n15327) );
NAND2_X1 U27682 ( .A1(n1452), .A2(n16070), .ZN(n1481) );
NAND2_X1 U27683 ( .A1(n16465), .A2(data_rdata_i_19_), .ZN(n1480) );
NAND2_X1 U27684 ( .A1(n1482), .A2(n1483), .ZN(n15326) );
NAND2_X1 U27685 ( .A1(n1452), .A2(n16071), .ZN(n1483) );
NAND2_X1 U27686 ( .A1(n16465), .A2(data_rdata_i_18_), .ZN(n1482) );
NAND2_X1 U27687 ( .A1(n1484), .A2(n1485), .ZN(n15325) );
NAND2_X1 U27688 ( .A1(n1452), .A2(n16072), .ZN(n1485) );
NAND2_X1 U27689 ( .A1(n16465), .A2(data_rdata_i_17_), .ZN(n1484) );
NAND2_X1 U27690 ( .A1(n1486), .A2(n1487), .ZN(n15324) );
NAND2_X1 U27691 ( .A1(n1452), .A2(n16073), .ZN(n1487) );
NAND2_X1 U27692 ( .A1(n16465), .A2(data_rdata_i_16_), .ZN(n1486) );
NAND2_X1 U27693 ( .A1(n1488), .A2(n1489), .ZN(n15323) );
NAND2_X1 U27694 ( .A1(n1452), .A2(n16074), .ZN(n1489) );
NAND2_X1 U27695 ( .A1(n16465), .A2(data_rdata_i_15_), .ZN(n1488) );
NAND2_X1 U27696 ( .A1(n1490), .A2(n1491), .ZN(n15322) );
NAND2_X1 U27697 ( .A1(n1452), .A2(n16075), .ZN(n1491) );
NAND2_X1 U27698 ( .A1(n16465), .A2(data_rdata_i_14_), .ZN(n1490) );
NAND2_X1 U27699 ( .A1(n1492), .A2(n1493), .ZN(n15321) );
NAND2_X1 U27700 ( .A1(n1452), .A2(n16076), .ZN(n1493) );
NAND2_X1 U27701 ( .A1(n16465), .A2(data_rdata_i_13_), .ZN(n1492) );
NAND2_X1 U27702 ( .A1(n1494), .A2(n1495), .ZN(n15320) );
NAND2_X1 U27703 ( .A1(n1452), .A2(n16077), .ZN(n1495) );
NAND2_X1 U27704 ( .A1(n16465), .A2(data_rdata_i_12_), .ZN(n1494) );
NAND2_X1 U27705 ( .A1(n1496), .A2(n1497), .ZN(n15319) );
NAND2_X1 U27706 ( .A1(n1452), .A2(n16078), .ZN(n1497) );
NAND2_X1 U27707 ( .A1(n16465), .A2(data_rdata_i_11_), .ZN(n1496) );
NAND2_X1 U27708 ( .A1(n1498), .A2(n1499), .ZN(n15318) );
NAND2_X1 U27709 ( .A1(n1452), .A2(n16079), .ZN(n1499) );
NAND2_X1 U27710 ( .A1(n16465), .A2(data_rdata_i_10_), .ZN(n1498) );
NAND2_X1 U27711 ( .A1(n1450), .A2(n1451), .ZN(n15317) );
NAND2_X1 U27712 ( .A1(n1452), .A2(n16080), .ZN(n1451) );
NAND2_X1 U27713 ( .A1(n16465), .A2(data_rdata_i_9_), .ZN(n1450) );
NAND2_X1 U27714 ( .A1(n7074), .A2(n7075), .ZN(n15772) );
NAND2_X1 U27715 ( .A1(n7072), .A2(n16195), .ZN(n7074) );
NAND2_X1 U27716 ( .A1(n19972), .A2(n6896), .ZN(n7075) );
NAND2_X1 U27717 ( .A1(n7070), .A2(n7071), .ZN(n14899) );
NAND2_X1 U27718 ( .A1(n7072), .A2(n16196), .ZN(n7070) );
NAND2_X1 U27719 ( .A1(n19972), .A2(n6943), .ZN(n7071) );
NAND2_X1 U27720 ( .A1(n5131), .A2(n5132), .ZN(n15557) );
NAND2_X1 U27721 ( .A1(n5133), .A2(n11498), .ZN(n5132) );
NAND2_X1 U27722 ( .A1(n7195), .A2(n7196), .ZN(n15394) );
OR2_X1 U27723 ( .A1(n7178), .A2(n11141), .ZN(n7196) );
NAND2_X1 U27724 ( .A1(n16397), .A2(n7037), .ZN(n7195) );
NAND2_X1 U27725 ( .A1(n7189), .A2(n7190), .ZN(n15393) );
OR2_X1 U27726 ( .A1(n16398), .A2(n11140), .ZN(n7190) );
NAND2_X1 U27727 ( .A1(n16397), .A2(n7191), .ZN(n7189) );
NAND2_X1 U27728 ( .A1(n7199), .A2(n7200), .ZN(n15388) );
OR2_X1 U27729 ( .A1(n16397), .A2(n11135), .ZN(n7200) );
NAND2_X1 U27730 ( .A1(n16397), .A2(n6803), .ZN(n7199) );
NAND2_X1 U27731 ( .A1(n7857), .A2(n7858), .ZN(n15361) );
OR2_X1 U27732 ( .A1(n16348), .A2(n11108), .ZN(n7858) );
NAND2_X1 U27733 ( .A1(n19977), .A2(n7068), .ZN(n7857) );
NAND2_X1 U27734 ( .A1(n7842), .A2(n7843), .ZN(n15114) );
OR2_X1 U27735 ( .A1(n19977), .A2(n10869), .ZN(n7843) );
NAND2_X1 U27736 ( .A1(n19977), .A2(n6925), .ZN(n7842) );
NAND2_X1 U27737 ( .A1(n7849), .A2(n7850), .ZN(n15082) );
OR2_X1 U27738 ( .A1(n19977), .A2(n10837), .ZN(n7850) );
NAND2_X1 U27739 ( .A1(n19977), .A2(n6952), .ZN(n7849) );
NAND2_X1 U27740 ( .A1(n7851), .A2(n7852), .ZN(n15068) );
OR2_X1 U27741 ( .A1(n16349), .A2(n10823), .ZN(n7852) );
NAND2_X1 U27742 ( .A1(n19977), .A2(n7237), .ZN(n7851) );
NAND2_X1 U27743 ( .A1(n7853), .A2(n7854), .ZN(n15053) );
OR2_X1 U27744 ( .A1(n16348), .A2(n10808), .ZN(n7854) );
NAND2_X1 U27745 ( .A1(n19977), .A2(n7240), .ZN(n7853) );
NAND2_X1 U27746 ( .A1(n7855), .A2(n7856), .ZN(n15039) );
OR2_X1 U27747 ( .A1(n19977), .A2(n10794), .ZN(n7856) );
NAND2_X1 U27748 ( .A1(n19977), .A2(n7243), .ZN(n7855) );
NAND2_X1 U27749 ( .A1(n7862), .A2(n7863), .ZN(n15000) );
OR2_X1 U27750 ( .A1(n19977), .A2(n10756), .ZN(n7863) );
NAND2_X1 U27751 ( .A1(n19977), .A2(n7250), .ZN(n7862) );
NAND2_X1 U27752 ( .A1(n7176), .A2(n7177), .ZN(n14987) );
OR2_X1 U27753 ( .A1(n16398), .A2(n10743), .ZN(n7177) );
NAND2_X1 U27754 ( .A1(n16397), .A2(n7179), .ZN(n7176) );
NAND2_X1 U27755 ( .A1(n7180), .A2(n7181), .ZN(n14973) );
OR2_X1 U27756 ( .A1(n16398), .A2(n10729), .ZN(n7181) );
NAND2_X1 U27757 ( .A1(n16397), .A2(n7182), .ZN(n7180) );
NAND2_X1 U27758 ( .A1(n7186), .A2(n7187), .ZN(n14959) );
OR2_X1 U27759 ( .A1(n7178), .A2(n10715), .ZN(n7187) );
NAND2_X1 U27760 ( .A1(n16397), .A2(n7188), .ZN(n7186) );
NAND2_X1 U27761 ( .A1(n7192), .A2(n7193), .ZN(n14946) );
OR2_X1 U27762 ( .A1(n16398), .A2(n10702), .ZN(n7193) );
NAND2_X1 U27763 ( .A1(n16397), .A2(n7194), .ZN(n7192) );
NAND2_X1 U27764 ( .A1(n7183), .A2(n7184), .ZN(n14934) );
OR2_X1 U27765 ( .A1(n7178), .A2(n10690), .ZN(n7184) );
NAND2_X1 U27766 ( .A1(n16397), .A2(n7185), .ZN(n7183) );
OR2_X1 U27767 ( .A1(n16274), .A2(n16275), .ZN(n15225) );
NOR2_X1 U27768 ( .A1(n7023), .A2(n10981), .ZN(n16274) );
NOR2_X1 U27769 ( .A1(n16400), .A2(n10980), .ZN(n16275) );
OR2_X1 U27770 ( .A1(n16276), .A2(n16277), .ZN(n15197) );
NOR2_X1 U27771 ( .A1(n7023), .A2(n10953), .ZN(n16276) );
NOR2_X1 U27772 ( .A1(n16400), .A2(n10952), .ZN(n16277) );
OR2_X1 U27773 ( .A1(n16278), .A2(n16279), .ZN(n15167) );
NOR2_X1 U27774 ( .A1(n7023), .A2(n10923), .ZN(n16278) );
NOR2_X1 U27775 ( .A1(n16400), .A2(n10922), .ZN(n16279) );
OR2_X1 U27776 ( .A1(n16280), .A2(n16281), .ZN(n15152) );
NOR2_X1 U27777 ( .A1(n7023), .A2(n10908), .ZN(n16280) );
NOR2_X1 U27778 ( .A1(n16400), .A2(n10907), .ZN(n16281) );
OR2_X1 U27779 ( .A1(n16282), .A2(n16283), .ZN(n14982) );
NOR2_X1 U27780 ( .A1(n7023), .A2(n10739), .ZN(n16282) );
NOR2_X1 U27781 ( .A1(n16400), .A2(n10738), .ZN(n16283) );
OR2_X1 U27782 ( .A1(n16284), .A2(n16285), .ZN(n14968) );
NOR2_X1 U27783 ( .A1(n7023), .A2(n10725), .ZN(n16284) );
NOR2_X1 U27784 ( .A1(n16400), .A2(n10724), .ZN(n16285) );
OR2_X1 U27785 ( .A1(n16286), .A2(n16287), .ZN(n14954) );
NOR2_X1 U27786 ( .A1(n16399), .A2(n10711), .ZN(n16286) );
NOR2_X1 U27787 ( .A1(n16400), .A2(n10710), .ZN(n16287) );
OR2_X1 U27788 ( .A1(n16288), .A2(n16289), .ZN(n14941) );
NOR2_X1 U27789 ( .A1(n7023), .A2(n10698), .ZN(n16288) );
NOR2_X1 U27790 ( .A1(n16401), .A2(n10697), .ZN(n16289) );
OR2_X1 U27791 ( .A1(n16290), .A2(n16291), .ZN(n14922) );
NOR2_X1 U27792 ( .A1(n7023), .A2(n10679), .ZN(n16290) );
NOR2_X1 U27793 ( .A1(n16400), .A2(n10678), .ZN(n16291) );
OR2_X1 U27794 ( .A1(n16292), .A2(n16293), .ZN(n14912) );
NOR2_X1 U27795 ( .A1(n16399), .A2(n10669), .ZN(n16292) );
NOR2_X1 U27796 ( .A1(n16401), .A2(n10668), .ZN(n16293) );
OR2_X1 U27797 ( .A1(n16294), .A2(n16295), .ZN(n14904) );
NOR2_X1 U27798 ( .A1(n7023), .A2(n10661), .ZN(n16294) );
NOR2_X1 U27799 ( .A1(n16400), .A2(n10660), .ZN(n16295) );
OR2_X1 U27800 ( .A1(n16296), .A2(n16297), .ZN(n14863) );
NOR2_X1 U27801 ( .A1(n7023), .A2(n10621), .ZN(n16296) );
NOR2_X1 U27802 ( .A1(n16401), .A2(n10620), .ZN(n16297) );
OR2_X1 U27803 ( .A1(n16298), .A2(n16299), .ZN(n14857) );
NOR2_X1 U27804 ( .A1(n7023), .A2(n10615), .ZN(n16298) );
NOR2_X1 U27805 ( .A1(n16400), .A2(n10614), .ZN(n16299) );
OR2_X1 U27806 ( .A1(n16300), .A2(n16301), .ZN(n14852) );
NOR2_X1 U27807 ( .A1(n7023), .A2(n10610), .ZN(n16300) );
NOR2_X1 U27808 ( .A1(n16401), .A2(n10609), .ZN(n16301) );
NAND2_X1 U27809 ( .A1(n6682), .A2(n6683), .ZN(n15268) );
OR2_X1 U27810 ( .A1(n6561), .A2(n11018), .ZN(n6683) );
NOR2_X1 U27811 ( .A1(n6684), .A2(n6685), .ZN(n6682) );
NOR2_X1 U27812 ( .A1(n19789), .A2(n6554), .ZN(n6684) );
NAND2_X1 U27813 ( .A1(n6586), .A2(n6587), .ZN(n15216) );
OR2_X1 U27814 ( .A1(n6561), .A2(n10971), .ZN(n6587) );
NOR2_X1 U27815 ( .A1(n6588), .A2(n6589), .ZN(n6586) );
NOR2_X1 U27816 ( .A1(n19757), .A2(n6554), .ZN(n6588) );
NAND2_X1 U27817 ( .A1(n6598), .A2(n6599), .ZN(n15186) );
OR2_X1 U27818 ( .A1(n6561), .A2(n10941), .ZN(n6599) );
NOR2_X1 U27819 ( .A1(n6600), .A2(n6601), .ZN(n6598) );
NOR2_X1 U27820 ( .A1(n19761), .A2(n6554), .ZN(n6600) );
NAND2_X1 U27821 ( .A1(n6628), .A2(n6629), .ZN(n15126) );
OR2_X1 U27822 ( .A1(n6561), .A2(n10881), .ZN(n6629) );
NOR2_X1 U27823 ( .A1(n6630), .A2(n6631), .ZN(n6628) );
NOR2_X1 U27824 ( .A1(n19771), .A2(n6554), .ZN(n6630) );
NAND2_X1 U27825 ( .A1(n6652), .A2(n6653), .ZN(n15079) );
OR2_X1 U27826 ( .A1(n6561), .A2(n10834), .ZN(n6653) );
NOR2_X1 U27827 ( .A1(n6654), .A2(n6655), .ZN(n6652) );
NOR2_X1 U27828 ( .A1(n19779), .A2(n6554), .ZN(n6654) );
NAND2_X1 U27829 ( .A1(n6580), .A2(n6581), .ZN(n14881) );
OR2_X1 U27830 ( .A1(n6561), .A2(n10638), .ZN(n6581) );
NOR2_X1 U27831 ( .A1(n6582), .A2(n6583), .ZN(n6580) );
NOR2_X1 U27832 ( .A1(n19755), .A2(n6554), .ZN(n6582) );
OR2_X1 U27833 ( .A1(n16302), .A2(n16303), .ZN(n15264) );
NOR2_X1 U27834 ( .A1(n16399), .A2(n11305), .ZN(n16302) );
NOR2_X1 U27835 ( .A1(n16401), .A2(n11304), .ZN(n16303) );
OR2_X1 U27836 ( .A1(n16304), .A2(n16305), .ZN(n15137) );
NOR2_X1 U27837 ( .A1(n16399), .A2(n10893), .ZN(n16304) );
NOR2_X1 U27838 ( .A1(n16401), .A2(n10892), .ZN(n16305) );
OR2_X1 U27839 ( .A1(n16306), .A2(n16307), .ZN(n15107) );
NOR2_X1 U27840 ( .A1(n16399), .A2(n10863), .ZN(n16306) );
NOR2_X1 U27841 ( .A1(n16401), .A2(n10862), .ZN(n16307) );
OR2_X1 U27842 ( .A1(n16308), .A2(n16309), .ZN(n15090) );
NOR2_X1 U27843 ( .A1(n7023), .A2(n10846), .ZN(n16308) );
NOR2_X1 U27844 ( .A1(n16401), .A2(n10845), .ZN(n16309) );
OR2_X1 U27845 ( .A1(n16310), .A2(n16311), .ZN(n15060) );
NOR2_X1 U27846 ( .A1(n16399), .A2(n10816), .ZN(n16310) );
NOR2_X1 U27847 ( .A1(n16401), .A2(n10815), .ZN(n16311) );
OR2_X1 U27848 ( .A1(n16312), .A2(n16313), .ZN(n15046) );
NOR2_X1 U27849 ( .A1(n16399), .A2(n10802), .ZN(n16312) );
NOR2_X1 U27850 ( .A1(n16401), .A2(n10801), .ZN(n16313) );
OR2_X1 U27851 ( .A1(n16314), .A2(n16315), .ZN(n15031) );
NOR2_X1 U27852 ( .A1(n16399), .A2(n10787), .ZN(n16314) );
NOR2_X1 U27853 ( .A1(n16401), .A2(n10786), .ZN(n16315) );
OR2_X1 U27854 ( .A1(n16316), .A2(n16317), .ZN(n15022) );
NOR2_X1 U27855 ( .A1(n16399), .A2(n10779), .ZN(n16316) );
NOR2_X1 U27856 ( .A1(n16401), .A2(n10778), .ZN(n16317) );
OR2_X1 U27857 ( .A1(n16318), .A2(n16319), .ZN(n15010) );
NOR2_X1 U27858 ( .A1(n16399), .A2(n10768), .ZN(n16318) );
NOR2_X1 U27859 ( .A1(n16401), .A2(n10767), .ZN(n16319) );
OR2_X1 U27860 ( .A1(n16320), .A2(n16321), .ZN(n14996) );
NOR2_X1 U27861 ( .A1(n16399), .A2(n10753), .ZN(n16320) );
NOR2_X1 U27862 ( .A1(n16401), .A2(n10752), .ZN(n16321) );
OR2_X1 U27863 ( .A1(n16322), .A2(n16323), .ZN(n14889) );
NOR2_X1 U27864 ( .A1(n7023), .A2(n10646), .ZN(n16322) );
NOR2_X1 U27865 ( .A1(n16401), .A2(n10645), .ZN(n16323) );
OR2_X1 U27866 ( .A1(n16324), .A2(n16325), .ZN(n14886) );
NOR2_X1 U27867 ( .A1(n16399), .A2(n10644), .ZN(n16324) );
NOR2_X1 U27868 ( .A1(n16401), .A2(n10643), .ZN(n16325) );
OR2_X1 U27869 ( .A1(n16326), .A2(n16327), .ZN(n14859) );
NOR2_X1 U27870 ( .A1(n7023), .A2(n10617), .ZN(n16326) );
NOR2_X1 U27871 ( .A1(n16401), .A2(n10616), .ZN(n16327) );
NAND2_X1 U27872 ( .A1(n7034), .A2(n7035), .ZN(n15754) );
NAND2_X1 U27873 ( .A1(n19972), .A2(n7037), .ZN(n7035) );
NOR2_X1 U27874 ( .A1(n7038), .A2(n7039), .ZN(n7034) );
NOR2_X1 U27875 ( .A1(n11477), .A2(n7040), .ZN(n7039) );
NAND2_X1 U27876 ( .A1(n3257), .A2(n3258), .ZN(n15641) );
OR2_X1 U27877 ( .A1(n19874), .A2(n11363), .ZN(n3258) );
NOR2_X1 U27878 ( .A1(n3260), .A2(n3261), .ZN(n3257) );
NOR2_X1 U27879 ( .A1(n19952), .A2(n3262), .ZN(n3261) );
NAND2_X1 U27880 ( .A1(n3264), .A2(n3265), .ZN(n15639) );
OR2_X1 U27881 ( .A1(n19874), .A2(n11361), .ZN(n3265) );
NOR2_X1 U27882 ( .A1(n3266), .A2(n3267), .ZN(n3264) );
NOR2_X1 U27883 ( .A1(n19953), .A2(n3262), .ZN(n3267) );
NAND2_X1 U27884 ( .A1(n3268), .A2(n3269), .ZN(n15637) );
OR2_X1 U27885 ( .A1(n19874), .A2(n11359), .ZN(n3269) );
NOR2_X1 U27886 ( .A1(n3270), .A2(n3271), .ZN(n3268) );
NOR2_X1 U27887 ( .A1(n19954), .A2(n3262), .ZN(n3271) );
NAND2_X1 U27888 ( .A1(n3272), .A2(n3273), .ZN(n15635) );
OR2_X1 U27889 ( .A1(n19874), .A2(n11357), .ZN(n3273) );
NOR2_X1 U27890 ( .A1(n3274), .A2(n3275), .ZN(n3272) );
NOR2_X1 U27891 ( .A1(n19955), .A2(n3262), .ZN(n3275) );
NAND2_X1 U27892 ( .A1(n3276), .A2(n3277), .ZN(n15633) );
OR2_X1 U27893 ( .A1(n19874), .A2(n11355), .ZN(n3277) );
NOR2_X1 U27894 ( .A1(n3278), .A2(n3279), .ZN(n3276) );
NOR2_X1 U27895 ( .A1(n19956), .A2(n3262), .ZN(n3279) );
NAND2_X1 U27896 ( .A1(n3280), .A2(n3281), .ZN(n15631) );
OR2_X1 U27897 ( .A1(n19874), .A2(n11353), .ZN(n3281) );
NOR2_X1 U27898 ( .A1(n3282), .A2(n3283), .ZN(n3280) );
NOR2_X1 U27899 ( .A1(n19957), .A2(n3262), .ZN(n3283) );
NAND2_X1 U27900 ( .A1(n3284), .A2(n3285), .ZN(n15629) );
OR2_X1 U27901 ( .A1(n19874), .A2(n11351), .ZN(n3285) );
NOR2_X1 U27902 ( .A1(n3286), .A2(n3287), .ZN(n3284) );
NOR2_X1 U27903 ( .A1(n19958), .A2(n3262), .ZN(n3287) );
NAND2_X1 U27904 ( .A1(n3297), .A2(n3298), .ZN(n15627) );
OR2_X1 U27905 ( .A1(n19874), .A2(n11349), .ZN(n3298) );
NOR2_X1 U27906 ( .A1(n3299), .A2(n3300), .ZN(n3297) );
NOR2_X1 U27907 ( .A1(n19959), .A2(n3262), .ZN(n3300) );
NAND2_X1 U27908 ( .A1(n2373), .A2(n2374), .ZN(n15575) );
NAND2_X1 U27909 ( .A1(rf_waddr_wb_o_4_), .A2(n16455), .ZN(n2373) );
NAND2_X1 U27910 ( .A1(n2375), .A2(n2103), .ZN(n2374) );
NAND2_X1 U27911 ( .A1(n2009), .A2(n2376), .ZN(n2375) );
NAND2_X1 U27912 ( .A1(n2412), .A2(n2726), .ZN(n15619) );
OR2_X1 U27913 ( .A1(n16453), .A2(n11341), .ZN(n2726) );
NAND2_X1 U27914 ( .A1(n2081), .A2(n2541), .ZN(n15581) );
OR2_X1 U27915 ( .A1(n16450), .A2(n11314), .ZN(n2541) );
NAND2_X1 U27916 ( .A1(n8457), .A2(n8458), .ZN(n15777) );
OR2_X1 U27917 ( .A1(n8452), .A2(n11508), .ZN(n8458) );
NOR2_X1 U27918 ( .A1(n8459), .A2(n8460), .ZN(n8457) );
AND2_X1 U27919 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_62), .A2(n8455), .ZN(n8460) );
NAND2_X1 U27920 ( .A1(n8178), .A2(n8179), .ZN(n15766) );
OR2_X1 U27921 ( .A1(n8165), .A2(n11490), .ZN(n8179) );
NOR2_X1 U27922 ( .A1(n8180), .A2(n8181), .ZN(n8178) );
AND2_X1 U27923 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_60), .A2(n8168), .ZN(n8181) );
NAND2_X1 U27924 ( .A1(n8410), .A2(n8411), .ZN(n15757) );
OR2_X1 U27925 ( .A1(n19979), .A2(n11479), .ZN(n8411) );
NOR2_X1 U27926 ( .A1(n8412), .A2(n8413), .ZN(n8410) );
AND2_X1 U27927 ( .A1(n11479), .A2(n8149), .ZN(n8413) );
NAND2_X1 U27928 ( .A1(n8210), .A2(n8211), .ZN(n15384) );
OR2_X1 U27929 ( .A1(n8165), .A2(n11131), .ZN(n8211) );
NOR2_X1 U27930 ( .A1(n8212), .A2(n8213), .ZN(n8210) );
AND2_X1 U27931 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_53), .A2(n8168), .ZN(n8213) );
NAND2_X1 U27932 ( .A1(n8358), .A2(n8359), .ZN(n15376) );
OR2_X1 U27933 ( .A1(n19979), .A2(n11123), .ZN(n8359) );
NOR2_X1 U27934 ( .A1(n8360), .A2(n8361), .ZN(n8358) );
AND2_X1 U27935 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_21), .A2(n16382), .ZN(n8361) );
NAND2_X1 U27936 ( .A1(n8366), .A2(n8367), .ZN(n15375) );
OR2_X1 U27937 ( .A1(n19979), .A2(n11122), .ZN(n8367) );
NOR2_X1 U27938 ( .A1(n8368), .A2(n8369), .ZN(n8366) );
AND2_X1 U27939 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_1), .A2(n16382), .ZN(n8369) );
NAND2_X1 U27940 ( .A1(n8497), .A2(n8498), .ZN(n15373) );
OR2_X1 U27941 ( .A1(n8452), .A2(n11120), .ZN(n8498) );
NOR2_X1 U27942 ( .A1(n8499), .A2(n8500), .ZN(n8497) );
AND2_X1 U27943 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_53), .A2(n8455), .ZN(n8500) );
NAND2_X1 U27944 ( .A1(n9298), .A2(n9299), .ZN(n15367) );
OR2_X1 U27945 ( .A1(n19981), .A2(n11114), .ZN(n9299) );
NOR2_X1 U27946 ( .A1(n9300), .A2(n9301), .ZN(n9298) );
AND2_X1 U27947 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_21), .A2(n8436), .ZN(n9301) );
NAND2_X1 U27948 ( .A1(n8186), .A2(n8187), .ZN(n15211) );
OR2_X1 U27949 ( .A1(n8165), .A2(n10966), .ZN(n8187) );
NOR2_X1 U27950 ( .A1(n8188), .A2(n8189), .ZN(n8186) );
AND2_X1 U27951 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_59), .A2(n8168), .ZN(n8189) );
NAND2_X1 U27952 ( .A1(n8473), .A2(n8474), .ZN(n15209) );
OR2_X1 U27953 ( .A1(n8452), .A2(n10964), .ZN(n8474) );
NOR2_X1 U27954 ( .A1(n8475), .A2(n8476), .ZN(n8473) );
AND2_X1 U27955 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_59), .A2(n8455), .ZN(n8476) );
NAND2_X1 U27956 ( .A1(n8190), .A2(n8191), .ZN(n15196) );
OR2_X1 U27957 ( .A1(n8165), .A2(n10951), .ZN(n8191) );
NOR2_X1 U27958 ( .A1(n8192), .A2(n8193), .ZN(n8190) );
AND2_X1 U27959 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_58), .A2(n8168), .ZN(n8193) );
NAND2_X1 U27960 ( .A1(n8477), .A2(n8478), .ZN(n15194) );
OR2_X1 U27961 ( .A1(n8452), .A2(n10949), .ZN(n8478) );
NOR2_X1 U27962 ( .A1(n8479), .A2(n8480), .ZN(n8477) );
AND2_X1 U27963 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_58), .A2(n8455), .ZN(n8480) );
NAND2_X1 U27964 ( .A1(n8194), .A2(n8195), .ZN(n15181) );
OR2_X1 U27965 ( .A1(n8165), .A2(n10936), .ZN(n8195) );
NOR2_X1 U27966 ( .A1(n8196), .A2(n8197), .ZN(n8194) );
AND2_X1 U27967 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_57), .A2(n8168), .ZN(n8197) );
NAND2_X1 U27968 ( .A1(n8342), .A2(n8343), .ZN(n15180) );
OR2_X1 U27969 ( .A1(n19979), .A2(n10935), .ZN(n8343) );
NOR2_X1 U27970 ( .A1(n8344), .A2(n8345), .ZN(n8342) );
AND2_X1 U27971 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_25), .A2(n16382), .ZN(n8345) );
NAND2_X1 U27972 ( .A1(n8481), .A2(n8482), .ZN(n15179) );
OR2_X1 U27973 ( .A1(n8452), .A2(n10934), .ZN(n8482) );
NOR2_X1 U27974 ( .A1(n8483), .A2(n8484), .ZN(n8481) );
AND2_X1 U27975 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_57), .A2(n8455), .ZN(n8484) );
NAND2_X1 U27976 ( .A1(n9134), .A2(n9135), .ZN(n15178) );
OR2_X1 U27977 ( .A1(n19981), .A2(n10933), .ZN(n9135) );
NOR2_X1 U27978 ( .A1(n9136), .A2(n9137), .ZN(n9134) );
AND2_X1 U27979 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_25), .A2(n8436), .ZN(n9137) );
NAND2_X1 U27980 ( .A1(n8198), .A2(n8199), .ZN(n15166) );
OR2_X1 U27981 ( .A1(n8165), .A2(n10921), .ZN(n8199) );
NOR2_X1 U27982 ( .A1(n8200), .A2(n8201), .ZN(n8198) );
AND2_X1 U27983 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_56), .A2(n8168), .ZN(n8201) );
NAND2_X1 U27984 ( .A1(n8346), .A2(n8347), .ZN(n15165) );
OR2_X1 U27985 ( .A1(n19979), .A2(n10920), .ZN(n8347) );
NOR2_X1 U27986 ( .A1(n8348), .A2(n8349), .ZN(n8346) );
AND2_X1 U27987 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_24), .A2(n16382), .ZN(n8349) );
NAND2_X1 U27988 ( .A1(n8485), .A2(n8486), .ZN(n15164) );
OR2_X1 U27989 ( .A1(n8452), .A2(n10919), .ZN(n8486) );
NOR2_X1 U27990 ( .A1(n8487), .A2(n8488), .ZN(n8485) );
AND2_X1 U27991 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_56), .A2(n8455), .ZN(n8488) );
NAND2_X1 U27992 ( .A1(n9175), .A2(n9176), .ZN(n15163) );
OR2_X1 U27993 ( .A1(n19981), .A2(n10918), .ZN(n9176) );
NOR2_X1 U27994 ( .A1(n9177), .A2(n9178), .ZN(n9175) );
AND2_X1 U27995 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_24), .A2(n8436), .ZN(n9178) );
NAND2_X1 U27996 ( .A1(n8202), .A2(n8203), .ZN(n15151) );
OR2_X1 U27997 ( .A1(n8165), .A2(n10906), .ZN(n8203) );
NOR2_X1 U27998 ( .A1(n8204), .A2(n8205), .ZN(n8202) );
AND2_X1 U27999 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_55), .A2(n8168), .ZN(n8205) );
NAND2_X1 U28000 ( .A1(n8350), .A2(n8351), .ZN(n15150) );
OR2_X1 U28001 ( .A1(n19979), .A2(n10905), .ZN(n8351) );
NOR2_X1 U28002 ( .A1(n8352), .A2(n8353), .ZN(n8350) );
AND2_X1 U28003 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_23), .A2(n16382), .ZN(n8353) );
NAND2_X1 U28004 ( .A1(n8489), .A2(n8490), .ZN(n15149) );
OR2_X1 U28005 ( .A1(n8452), .A2(n10904), .ZN(n8490) );
NOR2_X1 U28006 ( .A1(n8491), .A2(n8492), .ZN(n8489) );
AND2_X1 U28007 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_55), .A2(n8455), .ZN(n8492) );
NAND2_X1 U28008 ( .A1(n9216), .A2(n9217), .ZN(n15148) );
OR2_X1 U28009 ( .A1(n19981), .A2(n10903), .ZN(n9217) );
NOR2_X1 U28010 ( .A1(n9218), .A2(n9219), .ZN(n9216) );
AND2_X1 U28011 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_23), .A2(n8436), .ZN(n9219) );
NAND2_X1 U28012 ( .A1(n8206), .A2(n8207), .ZN(n15136) );
OR2_X1 U28013 ( .A1(n8165), .A2(n10891), .ZN(n8207) );
NOR2_X1 U28014 ( .A1(n8208), .A2(n8209), .ZN(n8206) );
AND2_X1 U28015 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_54), .A2(n8168), .ZN(n8209) );
NAND2_X1 U28016 ( .A1(n8354), .A2(n8355), .ZN(n15135) );
OR2_X1 U28017 ( .A1(n19979), .A2(n10890), .ZN(n8355) );
NOR2_X1 U28018 ( .A1(n8356), .A2(n8357), .ZN(n8354) );
AND2_X1 U28019 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_22), .A2(n16382), .ZN(n8357) );
NAND2_X1 U28020 ( .A1(n8493), .A2(n8494), .ZN(n15134) );
OR2_X1 U28021 ( .A1(n8452), .A2(n10889), .ZN(n8494) );
NOR2_X1 U28022 ( .A1(n8495), .A2(n8496), .ZN(n8493) );
AND2_X1 U28023 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_54), .A2(n8455), .ZN(n8496) );
NAND2_X1 U28024 ( .A1(n9257), .A2(n9258), .ZN(n15133) );
OR2_X1 U28025 ( .A1(n19981), .A2(n10888), .ZN(n9258) );
NOR2_X1 U28026 ( .A1(n9259), .A2(n9260), .ZN(n9257) );
AND2_X1 U28027 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_22), .A2(n8436), .ZN(n9260) );
NAND2_X1 U28028 ( .A1(n8214), .A2(n8215), .ZN(n15121) );
OR2_X1 U28029 ( .A1(n8165), .A2(n10876), .ZN(n8215) );
NOR2_X1 U28030 ( .A1(n8216), .A2(n8217), .ZN(n8214) );
AND2_X1 U28031 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_52), .A2(n8168), .ZN(n8217) );
NAND2_X1 U28032 ( .A1(n8362), .A2(n8363), .ZN(n15120) );
OR2_X1 U28033 ( .A1(n19979), .A2(n10875), .ZN(n8363) );
NOR2_X1 U28034 ( .A1(n8364), .A2(n8365), .ZN(n8362) );
AND2_X1 U28035 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_20), .A2(n16382), .ZN(n8365) );
NAND2_X1 U28036 ( .A1(n8501), .A2(n8502), .ZN(n15119) );
OR2_X1 U28037 ( .A1(n8452), .A2(n10874), .ZN(n8502) );
NOR2_X1 U28038 ( .A1(n8503), .A2(n8504), .ZN(n8501) );
AND2_X1 U28039 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_52), .A2(n8455), .ZN(n8504) );
NAND2_X1 U28040 ( .A1(n9341), .A2(n9342), .ZN(n15118) );
OR2_X1 U28041 ( .A1(n19981), .A2(n10873), .ZN(n9342) );
NOR2_X1 U28042 ( .A1(n9343), .A2(n9344), .ZN(n9341) );
AND2_X1 U28043 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_20), .A2(n8436), .ZN(n9344) );
NAND2_X1 U28044 ( .A1(n8218), .A2(n8219), .ZN(n15106) );
OR2_X1 U28045 ( .A1(n8165), .A2(n10861), .ZN(n8219) );
NOR2_X1 U28046 ( .A1(n8220), .A2(n8221), .ZN(n8218) );
AND2_X1 U28047 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_51), .A2(n8168), .ZN(n8221) );
NAND2_X1 U28048 ( .A1(n8370), .A2(n8371), .ZN(n15105) );
OR2_X1 U28049 ( .A1(n19979), .A2(n10860), .ZN(n8371) );
NOR2_X1 U28050 ( .A1(n8372), .A2(n8373), .ZN(n8370) );
AND2_X1 U28051 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_19), .A2(n16382), .ZN(n8373) );
NAND2_X1 U28052 ( .A1(n8505), .A2(n8506), .ZN(n15104) );
OR2_X1 U28053 ( .A1(n8452), .A2(n10859), .ZN(n8506) );
NOR2_X1 U28054 ( .A1(n8507), .A2(n8508), .ZN(n8505) );
AND2_X1 U28055 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_51), .A2(n8455), .ZN(n8508) );
NAND2_X1 U28056 ( .A1(n9428), .A2(n9429), .ZN(n15103) );
OR2_X1 U28057 ( .A1(n19981), .A2(n10858), .ZN(n9429) );
NOR2_X1 U28058 ( .A1(n9430), .A2(n9431), .ZN(n9428) );
AND2_X1 U28059 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_19), .A2(n8436), .ZN(n9431) );
NAND2_X1 U28060 ( .A1(n8222), .A2(n8223), .ZN(n15089) );
OR2_X1 U28061 ( .A1(n8165), .A2(n10844), .ZN(n8223) );
NOR2_X1 U28062 ( .A1(n8224), .A2(n8225), .ZN(n8222) );
AND2_X1 U28063 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_50), .A2(n8168), .ZN(n8225) );
NAND2_X1 U28064 ( .A1(n8374), .A2(n8375), .ZN(n15088) );
OR2_X1 U28065 ( .A1(n19979), .A2(n10843), .ZN(n8375) );
NOR2_X1 U28066 ( .A1(n8376), .A2(n8377), .ZN(n8374) );
AND2_X1 U28067 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_18), .A2(n16382), .ZN(n8377) );
NAND2_X1 U28068 ( .A1(n8509), .A2(n8510), .ZN(n15087) );
OR2_X1 U28069 ( .A1(n8452), .A2(n10842), .ZN(n8510) );
NOR2_X1 U28070 ( .A1(n8511), .A2(n8512), .ZN(n8509) );
AND2_X1 U28071 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_50), .A2(n8455), .ZN(n8512) );
NAND2_X1 U28072 ( .A1(n9469), .A2(n9470), .ZN(n15086) );
OR2_X1 U28073 ( .A1(n19981), .A2(n10841), .ZN(n9470) );
NOR2_X1 U28074 ( .A1(n9471), .A2(n9472), .ZN(n9469) );
AND2_X1 U28075 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_18), .A2(n8436), .ZN(n9472) );
NAND2_X1 U28076 ( .A1(n8234), .A2(n8235), .ZN(n15074) );
OR2_X1 U28077 ( .A1(n8165), .A2(n10829), .ZN(n8235) );
NOR2_X1 U28078 ( .A1(n8236), .A2(n8237), .ZN(n8234) );
AND2_X1 U28079 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_48), .A2(n8168), .ZN(n8237) );
NAND2_X1 U28080 ( .A1(n8382), .A2(n8383), .ZN(n15073) );
OR2_X1 U28081 ( .A1(n19979), .A2(n10828), .ZN(n8383) );
NOR2_X1 U28082 ( .A1(n8384), .A2(n8385), .ZN(n8382) );
AND2_X1 U28083 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_16), .A2(n8149), .ZN(n8385) );
NAND2_X1 U28084 ( .A1(n8521), .A2(n8522), .ZN(n15072) );
OR2_X1 U28085 ( .A1(n8452), .A2(n10827), .ZN(n8522) );
NOR2_X1 U28086 ( .A1(n8523), .A2(n8524), .ZN(n8521) );
AND2_X1 U28087 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_48), .A2(n8455), .ZN(n8524) );
NAND2_X1 U28088 ( .A1(n9554), .A2(n9555), .ZN(n15071) );
OR2_X1 U28089 ( .A1(n19981), .A2(n10826), .ZN(n9555) );
NOR2_X1 U28090 ( .A1(n9556), .A2(n9557), .ZN(n9554) );
AND2_X1 U28091 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_16), .A2(n8436), .ZN(n9557) );
NAND2_X1 U28092 ( .A1(n8238), .A2(n8239), .ZN(n15059) );
OR2_X1 U28093 ( .A1(n8165), .A2(n10814), .ZN(n8239) );
NOR2_X1 U28094 ( .A1(n8240), .A2(n8241), .ZN(n8238) );
AND2_X1 U28095 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_47), .A2(n8168), .ZN(n8241) );
NAND2_X1 U28096 ( .A1(n8386), .A2(n8387), .ZN(n15058) );
OR2_X1 U28097 ( .A1(n19979), .A2(n10813), .ZN(n8387) );
NOR2_X1 U28098 ( .A1(n8388), .A2(n8389), .ZN(n8386) );
AND2_X1 U28099 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_15), .A2(n8149), .ZN(n8389) );
NAND2_X1 U28100 ( .A1(n8525), .A2(n8526), .ZN(n15057) );
OR2_X1 U28101 ( .A1(n8452), .A2(n10812), .ZN(n8526) );
NOR2_X1 U28102 ( .A1(n8527), .A2(n8528), .ZN(n8525) );
AND2_X1 U28103 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_47), .A2(n8455), .ZN(n8528) );
NAND2_X1 U28104 ( .A1(n9596), .A2(n9597), .ZN(n15056) );
OR2_X1 U28105 ( .A1(n19981), .A2(n10811), .ZN(n9597) );
NOR2_X1 U28106 ( .A1(n9598), .A2(n9599), .ZN(n9596) );
AND2_X1 U28107 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_15), .A2(n16379), .ZN(n9599) );
NAND2_X1 U28108 ( .A1(n8242), .A2(n8243), .ZN(n15045) );
OR2_X1 U28109 ( .A1(n8165), .A2(n10800), .ZN(n8243) );
NOR2_X1 U28110 ( .A1(n8244), .A2(n8245), .ZN(n8242) );
AND2_X1 U28111 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_46), .A2(n8168), .ZN(n8245) );
NAND2_X1 U28112 ( .A1(n8390), .A2(n8391), .ZN(n15044) );
OR2_X1 U28113 ( .A1(n19979), .A2(n10799), .ZN(n8391) );
NOR2_X1 U28114 ( .A1(n8392), .A2(n8393), .ZN(n8390) );
AND2_X1 U28115 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_14), .A2(n8149), .ZN(n8393) );
NAND2_X1 U28116 ( .A1(n8529), .A2(n8530), .ZN(n15043) );
OR2_X1 U28117 ( .A1(n8452), .A2(n10798), .ZN(n8530) );
NOR2_X1 U28118 ( .A1(n8531), .A2(n8532), .ZN(n8529) );
AND2_X1 U28119 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_46), .A2(n8455), .ZN(n8532) );
NAND2_X1 U28120 ( .A1(n9634), .A2(n9635), .ZN(n15042) );
OR2_X1 U28121 ( .A1(n19981), .A2(n10797), .ZN(n9635) );
NOR2_X1 U28122 ( .A1(n9636), .A2(n9637), .ZN(n9634) );
AND2_X1 U28123 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_14), .A2(n8436), .ZN(n9637) );
NAND2_X1 U28124 ( .A1(n8394), .A2(n8395), .ZN(n15029) );
OR2_X1 U28125 ( .A1(n19979), .A2(n10784), .ZN(n8395) );
NOR2_X1 U28126 ( .A1(n8396), .A2(n8397), .ZN(n8394) );
AND2_X1 U28127 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_13), .A2(n8149), .ZN(n8397) );
NAND2_X1 U28128 ( .A1(n9671), .A2(n9672), .ZN(n15027) );
OR2_X1 U28129 ( .A1(n19981), .A2(n10782), .ZN(n9672) );
NOR2_X1 U28130 ( .A1(n9673), .A2(n9674), .ZN(n9671) );
AND2_X1 U28131 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_13), .A2(n16379), .ZN(n9674) );
NAND2_X1 U28132 ( .A1(n8398), .A2(n8399), .ZN(n15017) );
OR2_X1 U28133 ( .A1(n19979), .A2(n10774), .ZN(n8399) );
NOR2_X1 U28134 ( .A1(n8400), .A2(n8401), .ZN(n8398) );
AND2_X1 U28135 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_12), .A2(n8149), .ZN(n8401) );
NAND2_X1 U28136 ( .A1(n9708), .A2(n9709), .ZN(n15015) );
OR2_X1 U28137 ( .A1(n19981), .A2(n10772), .ZN(n9709) );
NOR2_X1 U28138 ( .A1(n9710), .A2(n9711), .ZN(n9708) );
AND2_X1 U28139 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_12), .A2(n8436), .ZN(n9711) );
NAND2_X1 U28140 ( .A1(n8402), .A2(n8403), .ZN(n15007) );
OR2_X1 U28141 ( .A1(n19979), .A2(n10763), .ZN(n8403) );
NOR2_X1 U28142 ( .A1(n8404), .A2(n8405), .ZN(n8402) );
AND2_X1 U28143 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_11), .A2(n8149), .ZN(n8405) );
NAND2_X1 U28144 ( .A1(n9748), .A2(n9749), .ZN(n15005) );
OR2_X1 U28145 ( .A1(n19981), .A2(n10761), .ZN(n9749) );
NOR2_X1 U28146 ( .A1(n9750), .A2(n9751), .ZN(n9748) );
AND2_X1 U28147 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_11), .A2(n16379), .ZN(n9751) );
NAND2_X1 U28148 ( .A1(n8406), .A2(n8407), .ZN(n14993) );
OR2_X1 U28149 ( .A1(n19979), .A2(n10749), .ZN(n8407) );
NOR2_X1 U28150 ( .A1(n8408), .A2(n8409), .ZN(n8406) );
AND2_X1 U28151 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_10), .A2(n8149), .ZN(n8409) );
NAND2_X1 U28152 ( .A1(n9796), .A2(n9797), .ZN(n14991) );
OR2_X1 U28153 ( .A1(n19981), .A2(n10747), .ZN(n9797) );
NOR2_X1 U28154 ( .A1(n9798), .A2(n9799), .ZN(n9796) );
AND2_X1 U28155 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_10), .A2(n8436), .ZN(n9799) );
NAND2_X1 U28156 ( .A1(n9383), .A2(n9384), .ZN(n14910) );
OR2_X1 U28157 ( .A1(n19981), .A2(n10666), .ZN(n9384) );
NOR2_X1 U28158 ( .A1(n9385), .A2(n9386), .ZN(n9383) );
AND2_X1 U28159 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_1), .A2(n8436), .ZN(n9386) );
NAND2_X1 U28160 ( .A1(n9833), .A2(n9834), .ZN(n14909) );
OR2_X1 U28161 ( .A1(n19981), .A2(n10665), .ZN(n9834) );
NOR2_X1 U28162 ( .A1(n9835), .A2(n9836), .ZN(n9833) );
AND2_X1 U28163 ( .A1(n10665), .A2(n16379), .ZN(n9836) );
NAND2_X1 U28164 ( .A1(n8230), .A2(n8231), .ZN(n14897) );
OR2_X1 U28165 ( .A1(n8165), .A2(n10653), .ZN(n8231) );
NOR2_X1 U28166 ( .A1(n8232), .A2(n8233), .ZN(n8230) );
AND2_X1 U28167 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_49), .A2(n8168), .ZN(n8233) );
NAND2_X1 U28168 ( .A1(n8378), .A2(n8379), .ZN(n14896) );
OR2_X1 U28169 ( .A1(n19979), .A2(n10652), .ZN(n8379) );
NOR2_X1 U28170 ( .A1(n8380), .A2(n8381), .ZN(n8378) );
AND2_X1 U28171 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_17), .A2(n16382), .ZN(n8381) );
NAND2_X1 U28172 ( .A1(n8517), .A2(n8518), .ZN(n14895) );
OR2_X1 U28173 ( .A1(n8452), .A2(n10651), .ZN(n8518) );
NOR2_X1 U28174 ( .A1(n8519), .A2(n8520), .ZN(n8517) );
AND2_X1 U28175 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_49), .A2(n8455), .ZN(n8520) );
NAND2_X1 U28176 ( .A1(n9510), .A2(n9511), .ZN(n14894) );
OR2_X1 U28177 ( .A1(n19981), .A2(n10650), .ZN(n9511) );
NOR2_X1 U28178 ( .A1(n9512), .A2(n9513), .ZN(n9510) );
AND2_X1 U28179 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_17), .A2(n8436), .ZN(n9513) );
NAND2_X1 U28180 ( .A1(n8465), .A2(n8466), .ZN(n14879) );
OR2_X1 U28181 ( .A1(n8452), .A2(n10636), .ZN(n8466) );
NOR2_X1 U28182 ( .A1(n8467), .A2(n8468), .ZN(n8465) );
AND2_X1 U28183 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_60), .A2(n8455), .ZN(n8468) );
NAND2_X1 U28184 ( .A1(n8174), .A2(n8175), .ZN(n14872) );
OR2_X1 U28185 ( .A1(n8165), .A2(n10629), .ZN(n8175) );
NOR2_X1 U28186 ( .A1(n8176), .A2(n8177), .ZN(n8174) );
AND2_X1 U28187 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_61), .A2(n8168), .ZN(n8177) );
NAND2_X1 U28188 ( .A1(n8170), .A2(n8171), .ZN(n14871) );
OR2_X1 U28189 ( .A1(n8165), .A2(n10628), .ZN(n8171) );
NOR2_X1 U28190 ( .A1(n8172), .A2(n8173), .ZN(n8170) );
AND2_X1 U28191 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_62), .A2(n8168), .ZN(n8173) );
NAND2_X1 U28192 ( .A1(n8163), .A2(n8164), .ZN(n14870) );
OR2_X1 U28193 ( .A1(n8165), .A2(n10627), .ZN(n8164) );
NOR2_X1 U28194 ( .A1(n8166), .A2(n8167), .ZN(n8163) );
AND2_X1 U28195 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_63), .A2(n8168), .ZN(n8167) );
NAND2_X1 U28196 ( .A1(n8461), .A2(n8462), .ZN(n14869) );
OR2_X1 U28197 ( .A1(n8452), .A2(n10626), .ZN(n8462) );
NOR2_X1 U28198 ( .A1(n8463), .A2(n8464), .ZN(n8461) );
AND2_X1 U28199 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_61), .A2(n8455), .ZN(n8464) );
NAND2_X1 U28200 ( .A1(n8450), .A2(n8451), .ZN(n14856) );
OR2_X1 U28201 ( .A1(n8452), .A2(n10613), .ZN(n8451) );
NOR2_X1 U28202 ( .A1(n8453), .A2(n8454), .ZN(n8450) );
AND2_X1 U28203 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_63), .A2(n8455), .ZN(n8454) );
NAND2_X1 U28204 ( .A1(n8091), .A2(n8092), .ZN(n15036) );
OR2_X1 U28205 ( .A1(n19969), .A2(n10791), .ZN(n8091) );
NAND2_X1 U28206 ( .A1(n19978), .A2(n7243), .ZN(n8092) );
NAND2_X1 U28207 ( .A1(n3020), .A2(n3021), .ZN(n15751) );
OR2_X1 U28208 ( .A1(n19886), .A2(n11472), .ZN(n3021) );
NAND2_X1 U28209 ( .A1(n19886), .A2(n15920), .ZN(n3020) );
NAND2_X1 U28210 ( .A1(n1512), .A2(n1513), .ZN(n15548) );
OR2_X1 U28211 ( .A1(n1514), .A2(n11294), .ZN(n1512) );
NAND2_X1 U28212 ( .A1(n1514), .A2(n1515), .ZN(n1513) );
NOR2_X1 U28213 ( .A1(n1511), .A2(n1520), .ZN(n1514) );
NAND2_X1 U28214 ( .A1(n2757), .A2(n2758), .ZN(n15761) );
OR2_X1 U28215 ( .A1(n1885), .A2(n11484), .ZN(n2758) );
NOR2_X1 U28216 ( .A1(n2759), .A2(n2760), .ZN(n2757) );
NOR2_X1 U28217 ( .A1(n2761), .A2(n16455), .ZN(n2760) );
NAND2_X1 U28218 ( .A1(n2242), .A2(n2667), .ZN(n15621) );
OR2_X1 U28219 ( .A1(n1885), .A2(n11343), .ZN(n2667) );
NAND2_X1 U28220 ( .A1(n8888), .A2(n8889), .ZN(n15778) );
OR2_X1 U28221 ( .A1(n19981), .A2(n11510), .ZN(n8889) );
NOR2_X1 U28222 ( .A1(n8890), .A2(n8891), .ZN(n8888) );
AND2_X1 U28223 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_31), .A2(n16379), .ZN(n8891) );
NAND2_X1 U28224 ( .A1(n8326), .A2(n8327), .ZN(n15767) );
OR2_X1 U28225 ( .A1(n19979), .A2(n11491), .ZN(n8327) );
NOR2_X1 U28226 ( .A1(n8328), .A2(n8329), .ZN(n8326) );
AND2_X1 U28227 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_29), .A2(n8149), .ZN(n8329) );
NAND2_X1 U28228 ( .A1(n8641), .A2(n8642), .ZN(n15755) );
OR2_X1 U28229 ( .A1(n19981), .A2(n11478), .ZN(n8642) );
NOR2_X1 U28230 ( .A1(n8643), .A2(n8644), .ZN(n8641) );
AND2_X1 U28231 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_3), .A2(n16379), .ZN(n8644) );
NAND2_X1 U28232 ( .A1(n8182), .A2(n8183), .ZN(n15385) );
OR2_X1 U28233 ( .A1(n19979), .A2(n11132), .ZN(n8183) );
NOR2_X1 U28234 ( .A1(n8184), .A2(n8185), .ZN(n8182) );
AND2_X1 U28235 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_5), .A2(n8149), .ZN(n8185) );
NAND2_X1 U28236 ( .A1(n8282), .A2(n8283), .ZN(n15383) );
OR2_X1 U28237 ( .A1(n8165), .A2(n11130), .ZN(n8283) );
NOR2_X1 U28238 ( .A1(n8284), .A2(n8285), .ZN(n8282) );
AND2_X1 U28239 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_37), .A2(n8168), .ZN(n8285) );
NAND2_X1 U28240 ( .A1(n8294), .A2(n8295), .ZN(n15382) );
OR2_X1 U28241 ( .A1(n8165), .A2(n11129), .ZN(n8295) );
NOR2_X1 U28242 ( .A1(n8296), .A2(n8297), .ZN(n8294) );
AND2_X1 U28243 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_34), .A2(n8168), .ZN(n8297) );
NAND2_X1 U28244 ( .A1(n8298), .A2(n8299), .ZN(n15381) );
OR2_X1 U28245 ( .A1(n8165), .A2(n11128), .ZN(n8299) );
NOR2_X1 U28246 ( .A1(n8300), .A2(n8301), .ZN(n8298) );
AND2_X1 U28247 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_33), .A2(n8168), .ZN(n8301) );
NAND2_X1 U28248 ( .A1(n8302), .A2(n8303), .ZN(n15380) );
OR2_X1 U28249 ( .A1(n8165), .A2(n11127), .ZN(n8303) );
NOR2_X1 U28250 ( .A1(n8304), .A2(n8305), .ZN(n8302) );
AND2_X1 U28251 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_32), .A2(n8168), .ZN(n8305) );
NAND2_X1 U28252 ( .A1(n8314), .A2(n8315), .ZN(n15379) );
OR2_X1 U28253 ( .A1(n19979), .A2(n11126), .ZN(n8315) );
NOR2_X1 U28254 ( .A1(n8316), .A2(n8317), .ZN(n8314) );
AND2_X1 U28255 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_31), .A2(n8149), .ZN(n8317) );
NAND2_X1 U28256 ( .A1(n8318), .A2(n8319), .ZN(n15378) );
OR2_X1 U28257 ( .A1(n19979), .A2(n11125), .ZN(n8319) );
NOR2_X1 U28258 ( .A1(n8320), .A2(n8321), .ZN(n8318) );
AND2_X1 U28259 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_30), .A2(n16382), .ZN(n8321) );
NAND2_X1 U28260 ( .A1(n8322), .A2(n8323), .ZN(n15377) );
OR2_X1 U28261 ( .A1(n19979), .A2(n11124), .ZN(n8323) );
NOR2_X1 U28262 ( .A1(n8324), .A2(n8325), .ZN(n8322) );
AND2_X1 U28263 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_2), .A2(n8149), .ZN(n8325) );
NAND2_X1 U28264 ( .A1(n8469), .A2(n8470), .ZN(n15374) );
OR2_X1 U28265 ( .A1(n19981), .A2(n11121), .ZN(n8470) );
NOR2_X1 U28266 ( .A1(n8471), .A2(n8472), .ZN(n8469) );
AND2_X1 U28267 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_5), .A2(n16379), .ZN(n8472) );
NAND2_X1 U28268 ( .A1(n8730), .A2(n8731), .ZN(n15372) );
OR2_X1 U28269 ( .A1(n8452), .A2(n11119), .ZN(n8731) );
NOR2_X1 U28270 ( .A1(n8732), .A2(n8733), .ZN(n8730) );
AND2_X1 U28271 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_37), .A2(n8455), .ZN(n8733) );
NAND2_X1 U28272 ( .A1(n8871), .A2(n8872), .ZN(n15371) );
OR2_X1 U28273 ( .A1(n8452), .A2(n11118), .ZN(n8872) );
NOR2_X1 U28274 ( .A1(n8873), .A2(n8874), .ZN(n8871) );
AND2_X1 U28275 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_34), .A2(n8455), .ZN(n8874) );
NAND2_X1 U28276 ( .A1(n8875), .A2(n8876), .ZN(n15370) );
OR2_X1 U28277 ( .A1(n8452), .A2(n11117), .ZN(n8876) );
NOR2_X1 U28278 ( .A1(n8877), .A2(n8878), .ZN(n8875) );
AND2_X1 U28279 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_33), .A2(n8455), .ZN(n8878) );
NAND2_X1 U28280 ( .A1(n8879), .A2(n8880), .ZN(n15369) );
OR2_X1 U28281 ( .A1(n8452), .A2(n11116), .ZN(n8880) );
NOR2_X1 U28282 ( .A1(n8881), .A2(n8882), .ZN(n8879) );
AND2_X1 U28283 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_32), .A2(n8455), .ZN(n8882) );
NAND2_X1 U28284 ( .A1(n8923), .A2(n8924), .ZN(n15368) );
OR2_X1 U28285 ( .A1(n19981), .A2(n11115), .ZN(n8924) );
NOR2_X1 U28286 ( .A1(n8925), .A2(n8926), .ZN(n8923) );
AND2_X1 U28287 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_30), .A2(n16379), .ZN(n8926) );
NAND2_X1 U28288 ( .A1(n8334), .A2(n8335), .ZN(n15210) );
OR2_X1 U28289 ( .A1(n19979), .A2(n10965), .ZN(n8335) );
NOR2_X1 U28290 ( .A1(n8336), .A2(n8337), .ZN(n8334) );
AND2_X1 U28291 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_27), .A2(n16382), .ZN(n8337) );
NAND2_X1 U28292 ( .A1(n9052), .A2(n9053), .ZN(n15208) );
OR2_X1 U28293 ( .A1(n19981), .A2(n10963), .ZN(n9053) );
NOR2_X1 U28294 ( .A1(n9054), .A2(n9055), .ZN(n9052) );
AND2_X1 U28295 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_27), .A2(n16379), .ZN(n9055) );
NAND2_X1 U28296 ( .A1(n8338), .A2(n8339), .ZN(n15195) );
OR2_X1 U28297 ( .A1(n19979), .A2(n10950), .ZN(n8339) );
NOR2_X1 U28298 ( .A1(n8340), .A2(n8341), .ZN(n8338) );
AND2_X1 U28299 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_26), .A2(n16382), .ZN(n8341) );
NAND2_X1 U28300 ( .A1(n9093), .A2(n9094), .ZN(n15193) );
OR2_X1 U28301 ( .A1(n19981), .A2(n10948), .ZN(n9094) );
NOR2_X1 U28302 ( .A1(n9095), .A2(n9096), .ZN(n9093) );
AND2_X1 U28303 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_26), .A2(n8436), .ZN(n9096) );
NAND2_X1 U28304 ( .A1(n8246), .A2(n8247), .ZN(n15030) );
OR2_X1 U28305 ( .A1(n8165), .A2(n10785), .ZN(n8247) );
NOR2_X1 U28306 ( .A1(n8248), .A2(n8249), .ZN(n8246) );
AND2_X1 U28307 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_45), .A2(n8168), .ZN(n8249) );
NAND2_X1 U28308 ( .A1(n8533), .A2(n8534), .ZN(n15028) );
OR2_X1 U28309 ( .A1(n8452), .A2(n10783), .ZN(n8534) );
NOR2_X1 U28310 ( .A1(n8535), .A2(n8536), .ZN(n8533) );
AND2_X1 U28311 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_45), .A2(n8455), .ZN(n8536) );
NAND2_X1 U28312 ( .A1(n8250), .A2(n8251), .ZN(n15018) );
OR2_X1 U28313 ( .A1(n8165), .A2(n10775), .ZN(n8251) );
NOR2_X1 U28314 ( .A1(n8252), .A2(n8253), .ZN(n8250) );
AND2_X1 U28315 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_44), .A2(n8168), .ZN(n8253) );
NAND2_X1 U28316 ( .A1(n8537), .A2(n8538), .ZN(n15016) );
OR2_X1 U28317 ( .A1(n8452), .A2(n10773), .ZN(n8538) );
NOR2_X1 U28318 ( .A1(n8539), .A2(n8540), .ZN(n8537) );
AND2_X1 U28319 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_44), .A2(n8455), .ZN(n8540) );
NAND2_X1 U28320 ( .A1(n8254), .A2(n8255), .ZN(n15008) );
OR2_X1 U28321 ( .A1(n8165), .A2(n10764), .ZN(n8255) );
NOR2_X1 U28322 ( .A1(n8256), .A2(n8257), .ZN(n8254) );
AND2_X1 U28323 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_43), .A2(n8168), .ZN(n8257) );
NAND2_X1 U28324 ( .A1(n8541), .A2(n8542), .ZN(n15006) );
OR2_X1 U28325 ( .A1(n8452), .A2(n10762), .ZN(n8542) );
NOR2_X1 U28326 ( .A1(n8543), .A2(n8544), .ZN(n8541) );
AND2_X1 U28327 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_43), .A2(n8455), .ZN(n8544) );
NAND2_X1 U28328 ( .A1(n8258), .A2(n8259), .ZN(n14994) );
OR2_X1 U28329 ( .A1(n8165), .A2(n10750), .ZN(n8259) );
NOR2_X1 U28330 ( .A1(n8260), .A2(n8261), .ZN(n8258) );
AND2_X1 U28331 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_42), .A2(n8168), .ZN(n8261) );
NAND2_X1 U28332 ( .A1(n8545), .A2(n8546), .ZN(n14992) );
OR2_X1 U28333 ( .A1(n8452), .A2(n10748), .ZN(n8546) );
NOR2_X1 U28334 ( .A1(n8547), .A2(n8548), .ZN(n8545) );
AND2_X1 U28335 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_42), .A2(n8455), .ZN(n8548) );
NAND2_X1 U28336 ( .A1(n8144), .A2(n8145), .ZN(n14980) );
OR2_X1 U28337 ( .A1(n19979), .A2(n10736), .ZN(n8145) );
NOR2_X1 U28338 ( .A1(n8147), .A2(n8148), .ZN(n8144) );
AND2_X1 U28339 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_9), .A2(n16382), .ZN(n8148) );
NAND2_X1 U28340 ( .A1(n8262), .A2(n8263), .ZN(n14979) );
OR2_X1 U28341 ( .A1(n8165), .A2(n10735), .ZN(n8263) );
NOR2_X1 U28342 ( .A1(n8264), .A2(n8265), .ZN(n8262) );
AND2_X1 U28343 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_41), .A2(n8168), .ZN(n8265) );
NAND2_X1 U28344 ( .A1(n8431), .A2(n8432), .ZN(n14978) );
OR2_X1 U28345 ( .A1(n19981), .A2(n10734), .ZN(n8432) );
NOR2_X1 U28346 ( .A1(n8434), .A2(n8435), .ZN(n8431) );
AND2_X1 U28347 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_9), .A2(n16379), .ZN(n8435) );
NAND2_X1 U28348 ( .A1(n8549), .A2(n8550), .ZN(n14977) );
OR2_X1 U28349 ( .A1(n8452), .A2(n10733), .ZN(n8550) );
NOR2_X1 U28350 ( .A1(n8551), .A2(n8552), .ZN(n8549) );
AND2_X1 U28351 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_41), .A2(n8455), .ZN(n8552) );
NAND2_X1 U28352 ( .A1(n8151), .A2(n8152), .ZN(n14966) );
OR2_X1 U28353 ( .A1(n19979), .A2(n10722), .ZN(n8152) );
NOR2_X1 U28354 ( .A1(n8153), .A2(n8154), .ZN(n8151) );
AND2_X1 U28355 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_8), .A2(n8149), .ZN(n8154) );
NAND2_X1 U28356 ( .A1(n8266), .A2(n8267), .ZN(n14965) );
OR2_X1 U28357 ( .A1(n8165), .A2(n10721), .ZN(n8267) );
NOR2_X1 U28358 ( .A1(n8268), .A2(n8269), .ZN(n8266) );
AND2_X1 U28359 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_40), .A2(n8168), .ZN(n8269) );
NAND2_X1 U28360 ( .A1(n8438), .A2(n8439), .ZN(n14964) );
OR2_X1 U28361 ( .A1(n19981), .A2(n10720), .ZN(n8439) );
NOR2_X1 U28362 ( .A1(n8440), .A2(n8441), .ZN(n8438) );
AND2_X1 U28363 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_8), .A2(n16379), .ZN(n8441) );
NAND2_X1 U28364 ( .A1(n8602), .A2(n8603), .ZN(n14963) );
OR2_X1 U28365 ( .A1(n8452), .A2(n10719), .ZN(n8603) );
NOR2_X1 U28366 ( .A1(n8604), .A2(n8605), .ZN(n8602) );
AND2_X1 U28367 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_40), .A2(n8455), .ZN(n8605) );
NAND2_X1 U28368 ( .A1(n8159), .A2(n8160), .ZN(n14953) );
OR2_X1 U28369 ( .A1(n19979), .A2(n10709), .ZN(n8160) );
NOR2_X1 U28370 ( .A1(n8161), .A2(n8162), .ZN(n8159) );
AND2_X1 U28371 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_6), .A2(n16382), .ZN(n8162) );
NAND2_X1 U28372 ( .A1(n8278), .A2(n8279), .ZN(n14952) );
OR2_X1 U28373 ( .A1(n8165), .A2(n10708), .ZN(n8279) );
NOR2_X1 U28374 ( .A1(n8280), .A2(n8281), .ZN(n8278) );
AND2_X1 U28375 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_38), .A2(n8168), .ZN(n8281) );
NAND2_X1 U28376 ( .A1(n8446), .A2(n8447), .ZN(n14951) );
OR2_X1 U28377 ( .A1(n19981), .A2(n10707), .ZN(n8447) );
NOR2_X1 U28378 ( .A1(n8448), .A2(n8449), .ZN(n8446) );
AND2_X1 U28379 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_6), .A2(n16379), .ZN(n8449) );
NAND2_X1 U28380 ( .A1(n8693), .A2(n8694), .ZN(n14950) );
OR2_X1 U28381 ( .A1(n8452), .A2(n10706), .ZN(n8694) );
NOR2_X1 U28382 ( .A1(n8695), .A2(n8696), .ZN(n8693) );
AND2_X1 U28383 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_38), .A2(n8455), .ZN(n8696) );
NAND2_X1 U28384 ( .A1(n8226), .A2(n8227), .ZN(n14940) );
OR2_X1 U28385 ( .A1(n19979), .A2(n10696), .ZN(n8227) );
NOR2_X1 U28386 ( .A1(n8228), .A2(n8229), .ZN(n8226) );
AND2_X1 U28387 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_4), .A2(n8149), .ZN(n8229) );
NAND2_X1 U28388 ( .A1(n8286), .A2(n8287), .ZN(n14939) );
OR2_X1 U28389 ( .A1(n8165), .A2(n10695), .ZN(n8287) );
NOR2_X1 U28390 ( .A1(n8288), .A2(n8289), .ZN(n8286) );
AND2_X1 U28391 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_36), .A2(n8168), .ZN(n8289) );
NAND2_X1 U28392 ( .A1(n8513), .A2(n8514), .ZN(n14938) );
OR2_X1 U28393 ( .A1(n19981), .A2(n10694), .ZN(n8514) );
NOR2_X1 U28394 ( .A1(n8515), .A2(n8516), .ZN(n8513) );
AND2_X1 U28395 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_4), .A2(n16379), .ZN(n8516) );
NAND2_X1 U28396 ( .A1(n8774), .A2(n8775), .ZN(n14937) );
OR2_X1 U28397 ( .A1(n8452), .A2(n10693), .ZN(n8775) );
NOR2_X1 U28398 ( .A1(n8776), .A2(n8777), .ZN(n8774) );
AND2_X1 U28399 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_36), .A2(n8455), .ZN(n8777) );
NAND2_X1 U28400 ( .A1(n8155), .A2(n8156), .ZN(n14930) );
OR2_X1 U28401 ( .A1(n19979), .A2(n10686), .ZN(n8156) );
NOR2_X1 U28402 ( .A1(n8157), .A2(n8158), .ZN(n8155) );
AND2_X1 U28403 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_7), .A2(n16382), .ZN(n8158) );
NAND2_X1 U28404 ( .A1(n8274), .A2(n8275), .ZN(n14929) );
OR2_X1 U28405 ( .A1(n8165), .A2(n10685), .ZN(n8275) );
NOR2_X1 U28406 ( .A1(n8276), .A2(n8277), .ZN(n8274) );
AND2_X1 U28407 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_39), .A2(n8168), .ZN(n8277) );
NAND2_X1 U28408 ( .A1(n8442), .A2(n8443), .ZN(n14928) );
OR2_X1 U28409 ( .A1(n19981), .A2(n10684), .ZN(n8443) );
NOR2_X1 U28410 ( .A1(n8444), .A2(n8445), .ZN(n8442) );
AND2_X1 U28411 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_7), .A2(n16379), .ZN(n8445) );
NAND2_X1 U28412 ( .A1(n8645), .A2(n8646), .ZN(n14927) );
OR2_X1 U28413 ( .A1(n8452), .A2(n10683), .ZN(n8646) );
NOR2_X1 U28414 ( .A1(n8647), .A2(n8648), .ZN(n8645) );
AND2_X1 U28415 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_39), .A2(n8455), .ZN(n8648) );
NAND2_X1 U28416 ( .A1(n8270), .A2(n8271), .ZN(n14919) );
OR2_X1 U28417 ( .A1(n19979), .A2(n10675), .ZN(n8271) );
NOR2_X1 U28418 ( .A1(n8272), .A2(n8273), .ZN(n8270) );
AND2_X1 U28419 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_3), .A2(n8149), .ZN(n8273) );
NAND2_X1 U28420 ( .A1(n8290), .A2(n8291), .ZN(n14918) );
OR2_X1 U28421 ( .A1(n8165), .A2(n10674), .ZN(n8291) );
NOR2_X1 U28422 ( .A1(n8292), .A2(n8293), .ZN(n8290) );
AND2_X1 U28423 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_35), .A2(n8168), .ZN(n8293) );
NAND2_X1 U28424 ( .A1(n8820), .A2(n8821), .ZN(n14917) );
OR2_X1 U28425 ( .A1(n8452), .A2(n10673), .ZN(n8821) );
NOR2_X1 U28426 ( .A1(n8822), .A2(n8823), .ZN(n8820) );
AND2_X1 U28427 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_35), .A2(n8455), .ZN(n8823) );
NAND2_X1 U28428 ( .A1(n8966), .A2(n8967), .ZN(n14911) );
OR2_X1 U28429 ( .A1(n19981), .A2(n10667), .ZN(n8967) );
NOR2_X1 U28430 ( .A1(n8968), .A2(n8969), .ZN(n8966) );
AND2_X1 U28431 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_2), .A2(n16379), .ZN(n8969) );
NAND2_X1 U28432 ( .A1(n8330), .A2(n8331), .ZN(n14880) );
OR2_X1 U28433 ( .A1(n19979), .A2(n10637), .ZN(n8331) );
NOR2_X1 U28434 ( .A1(n8332), .A2(n8333), .ZN(n8330) );
AND2_X1 U28435 ( .A1(cs_registers_i_minstret_counter_i_counter_upd_28), .A2(n16382), .ZN(n8333) );
NAND2_X1 U28436 ( .A1(n9011), .A2(n9012), .ZN(n14878) );
OR2_X1 U28437 ( .A1(n19981), .A2(n10635), .ZN(n9012) );
NOR2_X1 U28438 ( .A1(n9013), .A2(n9014), .ZN(n9011) );
AND2_X1 U28439 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_28), .A2(n16379), .ZN(n9014) );
NAND2_X1 U28440 ( .A1(n8970), .A2(n8971), .ZN(n14868) );
OR2_X1 U28441 ( .A1(n19981), .A2(n10625), .ZN(n8971) );
NOR2_X1 U28442 ( .A1(n8972), .A2(n8973), .ZN(n8970) );
AND2_X1 U28443 ( .A1(cs_registers_i_mcycle_counter_i_counter_upd_29), .A2(n16379), .ZN(n8973) );
NAND2_X1 U28444 ( .A1(n3253), .A2(n3254), .ZN(n15705) );
OR2_X1 U28445 ( .A1(n19873), .A2(n11424), .ZN(n3254) );
NOR2_X1 U28446 ( .A1(n3255), .A2(n3256), .ZN(n3253) );
NOR2_X1 U28447 ( .A1(n19961), .A2(n3129), .ZN(n3256) );
NAND2_X1 U28448 ( .A1(n3557), .A2(n3558), .ZN(n15704) );
OR2_X1 U28449 ( .A1(n19873), .A2(n11423), .ZN(n3558) );
NOR2_X1 U28450 ( .A1(n3559), .A2(n3560), .ZN(n3557) );
NOR2_X1 U28451 ( .A1(n11456), .A2(n16435), .ZN(n3560) );
NAND2_X1 U28452 ( .A1(n3156), .A2(n3157), .ZN(n15703) );
OR2_X1 U28453 ( .A1(n19873), .A2(n11422), .ZN(n3157) );
NOR2_X1 U28454 ( .A1(n3158), .A2(n3159), .ZN(n3156) );
NOR2_X1 U28455 ( .A1(n19908), .A2(n16436), .ZN(n3159) );
NAND2_X1 U28456 ( .A1(n3160), .A2(n3161), .ZN(n15702) );
OR2_X1 U28457 ( .A1(n19873), .A2(n11421), .ZN(n3161) );
NOR2_X1 U28458 ( .A1(n3162), .A2(n3163), .ZN(n3160) );
NOR2_X1 U28459 ( .A1(n19911), .A2(n16436), .ZN(n3163) );
NAND2_X1 U28460 ( .A1(n3168), .A2(n3169), .ZN(n15701) );
OR2_X1 U28461 ( .A1(n19873), .A2(n11420), .ZN(n3169) );
NOR2_X1 U28462 ( .A1(n3170), .A2(n3171), .ZN(n3168) );
NOR2_X1 U28463 ( .A1(n19913), .A2(n16436), .ZN(n3171) );
NAND2_X1 U28464 ( .A1(n3172), .A2(n3173), .ZN(n15700) );
OR2_X1 U28465 ( .A1(n19873), .A2(n11419), .ZN(n3173) );
NOR2_X1 U28466 ( .A1(n3174), .A2(n3175), .ZN(n3172) );
NOR2_X1 U28467 ( .A1(n19915), .A2(n16436), .ZN(n3175) );
NAND2_X1 U28468 ( .A1(n3176), .A2(n3177), .ZN(n15699) );
OR2_X1 U28469 ( .A1(n19873), .A2(n11418), .ZN(n3177) );
NOR2_X1 U28470 ( .A1(n3178), .A2(n3179), .ZN(n3176) );
NOR2_X1 U28471 ( .A1(n19918), .A2(n3129), .ZN(n3179) );
NAND2_X1 U28472 ( .A1(n3180), .A2(n3181), .ZN(n15698) );
OR2_X1 U28473 ( .A1(n19873), .A2(n11417), .ZN(n3181) );
NOR2_X1 U28474 ( .A1(n3182), .A2(n3183), .ZN(n3180) );
NOR2_X1 U28475 ( .A1(n19920), .A2(n3129), .ZN(n3183) );
NAND2_X1 U28476 ( .A1(n3184), .A2(n3185), .ZN(n15697) );
OR2_X1 U28477 ( .A1(n19873), .A2(n11416), .ZN(n3185) );
NOR2_X1 U28478 ( .A1(n3186), .A2(n3187), .ZN(n3184) );
NOR2_X1 U28479 ( .A1(n19922), .A2(n16436), .ZN(n3187) );
NAND2_X1 U28480 ( .A1(n3188), .A2(n3189), .ZN(n15696) );
OR2_X1 U28481 ( .A1(n19873), .A2(n11415), .ZN(n3189) );
NOR2_X1 U28482 ( .A1(n3190), .A2(n3191), .ZN(n3188) );
NOR2_X1 U28483 ( .A1(n19924), .A2(n3129), .ZN(n3191) );
NAND2_X1 U28484 ( .A1(n3192), .A2(n3193), .ZN(n15695) );
OR2_X1 U28485 ( .A1(n19873), .A2(n11414), .ZN(n3193) );
NOR2_X1 U28486 ( .A1(n3194), .A2(n3195), .ZN(n3192) );
NOR2_X1 U28487 ( .A1(n19926), .A2(n16436), .ZN(n3195) );
NAND2_X1 U28488 ( .A1(n3196), .A2(n3197), .ZN(n15694) );
OR2_X1 U28489 ( .A1(n19873), .A2(n11413), .ZN(n3197) );
NOR2_X1 U28490 ( .A1(n3198), .A2(n3199), .ZN(n3196) );
NOR2_X1 U28491 ( .A1(n19928), .A2(n3129), .ZN(n3199) );
NAND2_X1 U28492 ( .A1(n3200), .A2(n3201), .ZN(n15693) );
OR2_X1 U28493 ( .A1(n19873), .A2(n11412), .ZN(n3201) );
NOR2_X1 U28494 ( .A1(n3202), .A2(n3203), .ZN(n3200) );
NOR2_X1 U28495 ( .A1(n19930), .A2(n16436), .ZN(n3203) );
NAND2_X1 U28496 ( .A1(n3204), .A2(n3205), .ZN(n15692) );
OR2_X1 U28497 ( .A1(n19873), .A2(n11411), .ZN(n3205) );
NOR2_X1 U28498 ( .A1(n3206), .A2(n3207), .ZN(n3204) );
NOR2_X1 U28499 ( .A1(n19932), .A2(n3129), .ZN(n3207) );
NAND2_X1 U28500 ( .A1(n3212), .A2(n3213), .ZN(n15691) );
OR2_X1 U28501 ( .A1(n19873), .A2(n11410), .ZN(n3213) );
NOR2_X1 U28502 ( .A1(n3214), .A2(n3215), .ZN(n3212) );
NOR2_X1 U28503 ( .A1(n19933), .A2(n16436), .ZN(n3215) );
NAND2_X1 U28504 ( .A1(n3216), .A2(n3217), .ZN(n15690) );
OR2_X1 U28505 ( .A1(n19873), .A2(n11409), .ZN(n3217) );
NOR2_X1 U28506 ( .A1(n3218), .A2(n3219), .ZN(n3216) );
NOR2_X1 U28507 ( .A1(n19935), .A2(n3129), .ZN(n3219) );
NAND2_X1 U28508 ( .A1(n3220), .A2(n3221), .ZN(n15689) );
OR2_X1 U28509 ( .A1(n19873), .A2(n11408), .ZN(n3221) );
NOR2_X1 U28510 ( .A1(n3222), .A2(n3223), .ZN(n3220) );
NOR2_X1 U28511 ( .A1(n19944), .A2(n16436), .ZN(n3223) );
NAND2_X1 U28512 ( .A1(n3225), .A2(n3226), .ZN(n15688) );
OR2_X1 U28513 ( .A1(n19873), .A2(n11407), .ZN(n3226) );
NOR2_X1 U28514 ( .A1(n3227), .A2(n3228), .ZN(n3225) );
NOR2_X1 U28515 ( .A1(n19945), .A2(n3129), .ZN(n3228) );
NAND2_X1 U28516 ( .A1(n3233), .A2(n3234), .ZN(n15686) );
OR2_X1 U28517 ( .A1(n19873), .A2(n11405), .ZN(n3234) );
NOR2_X1 U28518 ( .A1(n3235), .A2(n3236), .ZN(n3233) );
NOR2_X1 U28519 ( .A1(n19947), .A2(n3129), .ZN(n3236) );
NAND2_X1 U28520 ( .A1(n3237), .A2(n3238), .ZN(n15685) );
OR2_X1 U28521 ( .A1(n19873), .A2(n11404), .ZN(n3238) );
NOR2_X1 U28522 ( .A1(n3239), .A2(n3240), .ZN(n3237) );
NOR2_X1 U28523 ( .A1(n19948), .A2(n3129), .ZN(n3240) );
NAND2_X1 U28524 ( .A1(n3241), .A2(n3242), .ZN(n15684) );
OR2_X1 U28525 ( .A1(n19873), .A2(n11403), .ZN(n3242) );
NOR2_X1 U28526 ( .A1(n3243), .A2(n3244), .ZN(n3241) );
NOR2_X1 U28527 ( .A1(n19949), .A2(n3129), .ZN(n3244) );
NAND2_X1 U28528 ( .A1(n3245), .A2(n3246), .ZN(n15683) );
OR2_X1 U28529 ( .A1(n19873), .A2(n11402), .ZN(n3246) );
NOR2_X1 U28530 ( .A1(n3247), .A2(n3248), .ZN(n3245) );
NOR2_X1 U28531 ( .A1(n19950), .A2(n3129), .ZN(n3248) );
NAND2_X1 U28532 ( .A1(n3249), .A2(n3250), .ZN(n15682) );
OR2_X1 U28533 ( .A1(n19873), .A2(n11401), .ZN(n3250) );
NOR2_X1 U28534 ( .A1(n3251), .A2(n3252), .ZN(n3249) );
NOR2_X1 U28535 ( .A1(n19951), .A2(n3129), .ZN(n3252) );
NAND2_X1 U28536 ( .A1(n3135), .A2(n3136), .ZN(n15679) );
OR2_X1 U28537 ( .A1(n19873), .A2(n11398), .ZN(n3136) );
NOR2_X1 U28538 ( .A1(n3138), .A2(n3139), .ZN(n3135) );
NOR2_X1 U28539 ( .A1(n19954), .A2(n16436), .ZN(n3139) );
NAND2_X1 U28540 ( .A1(n3148), .A2(n3149), .ZN(n15676) );
OR2_X1 U28541 ( .A1(n19873), .A2(n11395), .ZN(n3149) );
NOR2_X1 U28542 ( .A1(n3150), .A2(n3151), .ZN(n3148) );
NOR2_X1 U28543 ( .A1(n19957), .A2(n16436), .ZN(n3151) );
NAND2_X1 U28544 ( .A1(n3164), .A2(n3165), .ZN(n15674) );
OR2_X1 U28545 ( .A1(n19873), .A2(n11393), .ZN(n3165) );
NOR2_X1 U28546 ( .A1(n3166), .A2(n3167), .ZN(n3164) );
NOR2_X1 U28547 ( .A1(n19959), .A2(n16436), .ZN(n3167) );
NAND2_X1 U28548 ( .A1(n3571), .A2(n3572), .ZN(n15671) );
OR2_X1 U28549 ( .A1(n19874), .A2(n11390), .ZN(n3572) );
NOR2_X1 U28550 ( .A1(n3573), .A2(n3574), .ZN(n3571) );
NOR2_X1 U28551 ( .A1(n11423), .A2(n3263), .ZN(n3574) );
NAND2_X1 U28552 ( .A1(n3301), .A2(n3302), .ZN(n15668) );
OR2_X1 U28553 ( .A1(n19874), .A2(n11387), .ZN(n3302) );
NOR2_X1 U28554 ( .A1(n3303), .A2(n3304), .ZN(n3301) );
NOR2_X1 U28555 ( .A1(n19913), .A2(n3262), .ZN(n3304) );
NAND2_X1 U28556 ( .A1(n3305), .A2(n3306), .ZN(n15667) );
OR2_X1 U28557 ( .A1(n19874), .A2(n11386), .ZN(n3306) );
NOR2_X1 U28558 ( .A1(n3307), .A2(n3308), .ZN(n3305) );
NOR2_X1 U28559 ( .A1(n19915), .A2(n3262), .ZN(n3308) );
NAND2_X1 U28560 ( .A1(n3309), .A2(n3310), .ZN(n15666) );
OR2_X1 U28561 ( .A1(n19874), .A2(n11385), .ZN(n3310) );
NOR2_X1 U28562 ( .A1(n3311), .A2(n3312), .ZN(n3309) );
NOR2_X1 U28563 ( .A1(n19918), .A2(n16434), .ZN(n3312) );
NAND2_X1 U28564 ( .A1(n3313), .A2(n3314), .ZN(n15665) );
OR2_X1 U28565 ( .A1(n19874), .A2(n11462), .ZN(n3314) );
NOR2_X1 U28566 ( .A1(n3315), .A2(n3316), .ZN(n3313) );
NOR2_X1 U28567 ( .A1(n19920), .A2(n16434), .ZN(n3316) );
NAND2_X1 U28568 ( .A1(n3317), .A2(n3318), .ZN(n15664) );
OR2_X1 U28569 ( .A1(n19874), .A2(n11384), .ZN(n3318) );
NOR2_X1 U28570 ( .A1(n3319), .A2(n3320), .ZN(n3317) );
NOR2_X1 U28571 ( .A1(n19922), .A2(n16434), .ZN(n3320) );
NAND2_X1 U28572 ( .A1(n3325), .A2(n3326), .ZN(n15662) );
OR2_X1 U28573 ( .A1(n19874), .A2(n11382), .ZN(n3326) );
NOR2_X1 U28574 ( .A1(n3327), .A2(n3328), .ZN(n3325) );
NOR2_X1 U28575 ( .A1(n19926), .A2(n16434), .ZN(n3328) );
NAND2_X1 U28576 ( .A1(n3329), .A2(n3330), .ZN(n15661) );
OR2_X1 U28577 ( .A1(n19874), .A2(n11381), .ZN(n3330) );
NOR2_X1 U28578 ( .A1(n3331), .A2(n3332), .ZN(n3329) );
NOR2_X1 U28579 ( .A1(n19928), .A2(n16434), .ZN(n3332) );
NAND2_X1 U28580 ( .A1(n3337), .A2(n3338), .ZN(n15659) );
OR2_X1 U28581 ( .A1(n19874), .A2(n11379), .ZN(n3338) );
NOR2_X1 U28582 ( .A1(n3339), .A2(n3340), .ZN(n3337) );
NOR2_X1 U28583 ( .A1(n19932), .A2(n16434), .ZN(n3340) );
NAND2_X1 U28584 ( .A1(n3345), .A2(n3346), .ZN(n15658) );
OR2_X1 U28585 ( .A1(n19874), .A2(n11378), .ZN(n3346) );
NOR2_X1 U28586 ( .A1(n3347), .A2(n3348), .ZN(n3345) );
NOR2_X1 U28587 ( .A1(n19933), .A2(n16434), .ZN(n3348) );
NAND2_X1 U28588 ( .A1(n3349), .A2(n3350), .ZN(n15657) );
OR2_X1 U28589 ( .A1(n19874), .A2(n11377), .ZN(n3350) );
NOR2_X1 U28590 ( .A1(n3351), .A2(n3352), .ZN(n3349) );
NOR2_X1 U28591 ( .A1(n19935), .A2(n16434), .ZN(n3352) );
NAND2_X1 U28592 ( .A1(n3363), .A2(n3364), .ZN(n15652) );
OR2_X1 U28593 ( .A1(n19874), .A2(n11373), .ZN(n3364) );
NOR2_X1 U28594 ( .A1(n3365), .A2(n3366), .ZN(n3363) );
NOR2_X1 U28595 ( .A1(n19946), .A2(n3262), .ZN(n3366) );
NAND2_X1 U28596 ( .A1(n3367), .A2(n3368), .ZN(n15650) );
OR2_X1 U28597 ( .A1(n19874), .A2(n11371), .ZN(n3368) );
NOR2_X1 U28598 ( .A1(n3369), .A2(n3370), .ZN(n3367) );
NOR2_X1 U28599 ( .A1(n19947), .A2(n16434), .ZN(n3370) );
NAND2_X1 U28600 ( .A1(n3371), .A2(n3372), .ZN(n15648) );
OR2_X1 U28601 ( .A1(n19874), .A2(n11369), .ZN(n3372) );
NOR2_X1 U28602 ( .A1(n3373), .A2(n3374), .ZN(n3371) );
NOR2_X1 U28603 ( .A1(n19948), .A2(n3262), .ZN(n3374) );
NAND2_X1 U28604 ( .A1(n3375), .A2(n3376), .ZN(n15646) );
OR2_X1 U28605 ( .A1(n19874), .A2(n11367), .ZN(n3376) );
NOR2_X1 U28606 ( .A1(n3377), .A2(n3378), .ZN(n3375) );
NOR2_X1 U28607 ( .A1(n19949), .A2(n16434), .ZN(n3378) );
NAND2_X1 U28608 ( .A1(n3379), .A2(n3380), .ZN(n15644) );
OR2_X1 U28609 ( .A1(n19874), .A2(n11365), .ZN(n3380) );
NOR2_X1 U28610 ( .A1(n3381), .A2(n3382), .ZN(n3379) );
NOR2_X1 U28611 ( .A1(n19950), .A2(n3262), .ZN(n3382) );
NAND2_X1 U28612 ( .A1(n3383), .A2(n3384), .ZN(n15642) );
OR2_X1 U28613 ( .A1(n19874), .A2(n11461), .ZN(n3384) );
NOR2_X1 U28614 ( .A1(n3385), .A2(n3386), .ZN(n3383) );
NOR2_X1 U28615 ( .A1(n19951), .A2(n16434), .ZN(n3386) );
NAND2_X1 U28616 ( .A1(n1529), .A2(n1530), .ZN(n15549) );
OR2_X1 U28617 ( .A1(n1531), .A2(n11295), .ZN(n1530) );
NAND2_X1 U28618 ( .A1(n1525), .A2(data_gnt_i), .ZN(n1529) );
NAND2_X1 U28619 ( .A1(n7747), .A2(n7748), .ZN(n15348) );
OR2_X1 U28620 ( .A1(n19976), .A2(n11095), .ZN(n7748) );
NAND2_X1 U28621 ( .A1(n16347), .A2(n6824), .ZN(n7747) );
NAND2_X1 U28622 ( .A1(n7743), .A2(n7744), .ZN(n15347) );
OR2_X1 U28623 ( .A1(n16347), .A2(n11094), .ZN(n7744) );
NAND2_X1 U28624 ( .A1(n16347), .A2(n6803), .ZN(n7743) );
NAND2_X1 U28625 ( .A1(n5117), .A2(n5118), .ZN(n15254) );
OR2_X1 U28626 ( .A1(n5119), .A2(n5120), .ZN(n5118) );
NAND2_X1 U28627 ( .A1(nmi_mode), .A2(n5119), .ZN(n5117) );
NAND2_X1 U28628 ( .A1(n5121), .A2(n5122), .ZN(n5119) );
NAND2_X1 U28629 ( .A1(n7567), .A2(n7568), .ZN(n15253) );
NAND2_X1 U28630 ( .A1(n15808), .A2(crash_dump_o_0_), .ZN(n7568) );
NOR2_X1 U28631 ( .A1(n7572), .A2(n7573), .ZN(n7567) );
NOR2_X1 U28632 ( .A1(n11464), .A2(n16392), .ZN(n7573) );
NAND2_X1 U28633 ( .A1(n1545), .A2(n1546), .ZN(n15552) );
NOR2_X1 U28634 ( .A1(n1551), .A2(n1552), .ZN(n1545) );
NOR2_X1 U28635 ( .A1(n1547), .A2(n1548), .ZN(n1546) );
NOR2_X1 U28636 ( .A1(data_gnt_i), .A2(n1541), .ZN(n1552) );
NAND2_X1 U28637 ( .A1(n1591), .A2(n1592), .ZN(n15316) );
OR2_X1 U28638 ( .A1(n19963), .A2(n11065), .ZN(n1591) );
NAND2_X1 U28639 ( .A1(n1593), .A2(n1594), .ZN(n1592) );
NOR2_X1 U28640 ( .A1(n15805), .A2(n1596), .ZN(n1594) );
NAND2_X1 U28641 ( .A1(n2197), .A2(n2198), .ZN(n15607) );
NOR2_X1 U28642 ( .A1(n2206), .A2(n2207), .ZN(n2197) );
NOR2_X1 U28643 ( .A1(n2178), .A2(n2199), .ZN(n2198) );
NOR2_X1 U28644 ( .A1(n11331), .A2(n16453), .ZN(n2207) );
NAND2_X1 U28645 ( .A1(n2732), .A2(n2733), .ZN(n14888) );
NAND2_X1 U28646 ( .A1(n16457), .A2(instr_fetch_err_plus2), .ZN(n2732) );
NAND2_X1 U28647 ( .A1(n2734), .A2(n11390), .ZN(n2733) );
NOR2_X1 U28648 ( .A1(n2735), .A2(n16457), .ZN(n2734) );
NAND2_X1 U28649 ( .A1(n7150), .A2(n7151), .ZN(n15263) );
OR2_X1 U28650 ( .A1(n16399), .A2(n11476), .ZN(n7150) );
NAND2_X1 U28651 ( .A1(n7023), .A2(n16081), .ZN(n7151) );
NAND2_X1 U28652 ( .A1(n2077), .A2(n2078), .ZN(n15590) );
NOR2_X1 U28653 ( .A1(n19878), .A2(n2080), .ZN(n2077) );
NOR2_X1 U28654 ( .A1(n11501), .A2(n16450), .ZN(n2080) );
NAND2_X1 U28655 ( .A1(n2533), .A2(n2078), .ZN(n15589) );
NOR2_X1 U28656 ( .A1(n19878), .A2(n2540), .ZN(n2533) );
NOR2_X1 U28657 ( .A1(n11321), .A2(n16450), .ZN(n2540) );
NAND2_X1 U28658 ( .A1(n8068), .A2(n8069), .ZN(n15228) );
OR2_X1 U28659 ( .A1(n20988), .A2(n10983), .ZN(n8068) );
NAND2_X1 U28660 ( .A1(n8070), .A2(n15909), .ZN(n8069) );
NAND2_X1 U28661 ( .A1(n8072), .A2(n8073), .ZN(n15227) );
OR2_X1 U28662 ( .A1(n20988), .A2(n10982), .ZN(n8072) );
NAND2_X1 U28663 ( .A1(n8070), .A2(n11301), .ZN(n8073) );
NAND2_X1 U28664 ( .A1(n2020), .A2(n2021), .ZN(n15618) );
NAND2_X1 U28665 ( .A1(rf_waddr_wb_o_1_), .A2(n16454), .ZN(n2021) );
NOR2_X1 U28666 ( .A1(n2022), .A2(n2023), .ZN(n2020) );
NOR2_X1 U28667 ( .A1(n2027), .A2(n2028), .ZN(n2022) );
NAND2_X1 U28668 ( .A1(n2031), .A2(n2032), .ZN(n15617) );
NAND2_X1 U28669 ( .A1(rf_waddr_wb_o_0_), .A2(n16457), .ZN(n2032) );
NOR2_X1 U28670 ( .A1(n2033), .A2(n2034), .ZN(n2031) );
NOR2_X1 U28671 ( .A1(n2037), .A2(n16456), .ZN(n2033) );
NAND2_X1 U28672 ( .A1(n2004), .A2(n2005), .ZN(n15576) );
NAND2_X1 U28673 ( .A1(rf_waddr_wb_o_2_), .A2(n16456), .ZN(n2005) );
NOR2_X1 U28674 ( .A1(n2006), .A2(n2007), .ZN(n2004) );
NOR2_X1 U28675 ( .A1(n19921), .A2(n2009), .ZN(n2007) );
NAND2_X1 U28676 ( .A1(n3711), .A2(n3712), .ZN(n15747) );
NOR2_X1 U28677 ( .A1(n3719), .A2(n3720), .ZN(n3711) );
NOR2_X1 U28678 ( .A1(n3713), .A2(n3714), .ZN(n3712) );
NOR2_X1 U28679 ( .A1(n11468), .A2(n3019), .ZN(n3720) );
NAND2_X1 U28680 ( .A1(n8045), .A2(n8046), .ZN(n15567) );
NOR2_X1 U28681 ( .A1(n8049), .A2(n8050), .ZN(n8045) );
NOR2_X1 U28682 ( .A1(n8047), .A2(n8048), .ZN(n8046) );
NOR2_X1 U28683 ( .A1(n11306), .A2(n7875), .ZN(n8050) );
NAND2_X1 U28684 ( .A1(n8015), .A2(n8016), .ZN(n15085) );
NOR2_X1 U28685 ( .A1(n8019), .A2(n8020), .ZN(n8015) );
NOR2_X1 U28686 ( .A1(n8017), .A2(n8018), .ZN(n8016) );
NOR2_X1 U28687 ( .A1(n10840), .A2(n16388), .ZN(n8020) );
NAND2_X1 U28688 ( .A1(n8021), .A2(n8022), .ZN(n15070) );
NOR2_X1 U28689 ( .A1(n8025), .A2(n8026), .ZN(n8021) );
NOR2_X1 U28690 ( .A1(n8023), .A2(n8024), .ZN(n8022) );
NOR2_X1 U28691 ( .A1(n10825), .A2(n7875), .ZN(n8026) );
NAND2_X1 U28692 ( .A1(n8027), .A2(n8028), .ZN(n15055) );
NOR2_X1 U28693 ( .A1(n8031), .A2(n8032), .ZN(n8027) );
NOR2_X1 U28694 ( .A1(n8029), .A2(n8030), .ZN(n8028) );
NOR2_X1 U28695 ( .A1(n10810), .A2(n16388), .ZN(n8032) );
NAND2_X1 U28696 ( .A1(n8033), .A2(n8034), .ZN(n15041) );
NOR2_X1 U28697 ( .A1(n8037), .A2(n8038), .ZN(n8033) );
NOR2_X1 U28698 ( .A1(n8035), .A2(n8036), .ZN(n8034) );
NOR2_X1 U28699 ( .A1(n10796), .A2(n7875), .ZN(n8038) );
NAND2_X1 U28700 ( .A1(n8039), .A2(n8040), .ZN(n15014) );
NOR2_X1 U28701 ( .A1(n8043), .A2(n8044), .ZN(n8039) );
NOR2_X1 U28702 ( .A1(n8041), .A2(n8042), .ZN(n8040) );
NOR2_X1 U28703 ( .A1(n10771), .A2(n16388), .ZN(n8044) );
NAND2_X1 U28704 ( .A1(n8051), .A2(n8052), .ZN(n15002) );
NOR2_X1 U28705 ( .A1(n8057), .A2(n8058), .ZN(n8051) );
NOR2_X1 U28706 ( .A1(n8053), .A2(n8054), .ZN(n8052) );
NOR2_X1 U28707 ( .A1(n10758), .A2(n7875), .ZN(n8058) );
NAND2_X1 U28708 ( .A1(n6818), .A2(n6819), .ZN(n15768) );
NOR2_X1 U28709 ( .A1(n6825), .A2(n6826), .ZN(n6818) );
NOR2_X1 U28710 ( .A1(n6820), .A2(n6821), .ZN(n6819) );
NOR2_X1 U28711 ( .A1(n11494), .A2(n6719), .ZN(n6826) );
NAND2_X1 U28712 ( .A1(n6890), .A2(n6891), .ZN(n15259) );
NOR2_X1 U28713 ( .A1(n6897), .A2(n6898), .ZN(n6890) );
NOR2_X1 U28714 ( .A1(n6892), .A2(n6893), .ZN(n6891) );
NOR2_X1 U28715 ( .A1(n11013), .A2(n16402), .ZN(n6898) );
NAND2_X1 U28716 ( .A1(n6836), .A2(n6837), .ZN(n15217) );
NOR2_X1 U28717 ( .A1(n6843), .A2(n6844), .ZN(n6836) );
NOR2_X1 U28718 ( .A1(n6838), .A2(n6839), .ZN(n6837) );
NOR2_X1 U28719 ( .A1(n10972), .A2(n6719), .ZN(n6844) );
NAND2_X1 U28720 ( .A1(n6845), .A2(n6846), .ZN(n15202) );
NOR2_X1 U28721 ( .A1(n6852), .A2(n6853), .ZN(n6845) );
NOR2_X1 U28722 ( .A1(n6847), .A2(n6848), .ZN(n6846) );
NOR2_X1 U28723 ( .A1(n10957), .A2(n16402), .ZN(n6853) );
NAND2_X1 U28724 ( .A1(n6854), .A2(n6855), .ZN(n15187) );
NOR2_X1 U28725 ( .A1(n6861), .A2(n6862), .ZN(n6854) );
NOR2_X1 U28726 ( .A1(n6856), .A2(n6857), .ZN(n6855) );
NOR2_X1 U28727 ( .A1(n10942), .A2(n6719), .ZN(n6862) );
NAND2_X1 U28728 ( .A1(n6863), .A2(n6864), .ZN(n15172) );
NOR2_X1 U28729 ( .A1(n6870), .A2(n6871), .ZN(n6863) );
NOR2_X1 U28730 ( .A1(n6865), .A2(n6866), .ZN(n6864) );
NOR2_X1 U28731 ( .A1(n10927), .A2(n16402), .ZN(n6871) );
NAND2_X1 U28732 ( .A1(n6872), .A2(n6873), .ZN(n15157) );
NOR2_X1 U28733 ( .A1(n6879), .A2(n6880), .ZN(n6872) );
NOR2_X1 U28734 ( .A1(n6874), .A2(n6875), .ZN(n6873) );
NOR2_X1 U28735 ( .A1(n10912), .A2(n6719), .ZN(n6880) );
NAND2_X1 U28736 ( .A1(n6881), .A2(n6882), .ZN(n15142) );
NOR2_X1 U28737 ( .A1(n6888), .A2(n6889), .ZN(n6881) );
NOR2_X1 U28738 ( .A1(n6883), .A2(n6884), .ZN(n6882) );
NOR2_X1 U28739 ( .A1(n10897), .A2(n16402), .ZN(n6889) );
NAND2_X1 U28740 ( .A1(n6899), .A2(n6900), .ZN(n15127) );
NOR2_X1 U28741 ( .A1(n6906), .A2(n6907), .ZN(n6899) );
NOR2_X1 U28742 ( .A1(n6901), .A2(n6902), .ZN(n6900) );
NOR2_X1 U28743 ( .A1(n10882), .A2(n6719), .ZN(n6907) );
NAND2_X1 U28744 ( .A1(n6919), .A2(n6920), .ZN(n15112) );
NOR2_X1 U28745 ( .A1(n6926), .A2(n6927), .ZN(n6919) );
NOR2_X1 U28746 ( .A1(n6921), .A2(n6922), .ZN(n6920) );
NOR2_X1 U28747 ( .A1(n10867), .A2(n16402), .ZN(n6927) );
NAND2_X1 U28748 ( .A1(n6928), .A2(n6929), .ZN(n15095) );
NOR2_X1 U28749 ( .A1(n6935), .A2(n6936), .ZN(n6928) );
NOR2_X1 U28750 ( .A1(n6930), .A2(n6931), .ZN(n6929) );
NOR2_X1 U28751 ( .A1(n10850), .A2(n16402), .ZN(n6936) );
NAND2_X1 U28752 ( .A1(n6946), .A2(n6947), .ZN(n15080) );
NOR2_X1 U28753 ( .A1(n6953), .A2(n6954), .ZN(n6946) );
NOR2_X1 U28754 ( .A1(n6948), .A2(n6949), .ZN(n6947) );
NOR2_X1 U28755 ( .A1(n10835), .A2(n16402), .ZN(n6954) );
NAND2_X1 U28756 ( .A1(n6937), .A2(n6938), .ZN(n14900) );
NOR2_X1 U28757 ( .A1(n6944), .A2(n6945), .ZN(n6937) );
NOR2_X1 U28758 ( .A1(n6939), .A2(n6940), .ZN(n6938) );
NOR2_X1 U28759 ( .A1(n10656), .A2(n16402), .ZN(n6945) );
NAND2_X1 U28760 ( .A1(n6827), .A2(n6828), .ZN(n14882) );
NOR2_X1 U28761 ( .A1(n6834), .A2(n6835), .ZN(n6827) );
NOR2_X1 U28762 ( .A1(n6829), .A2(n6830), .ZN(n6828) );
NOR2_X1 U28763 ( .A1(n10639), .A2(n16402), .ZN(n6835) );
NAND2_X1 U28764 ( .A1(n6797), .A2(n6798), .ZN(n14862) );
NOR2_X1 U28765 ( .A1(n6804), .A2(n6805), .ZN(n6797) );
NOR2_X1 U28766 ( .A1(n6799), .A2(n6800), .ZN(n6798) );
NOR2_X1 U28767 ( .A1(n10619), .A2(n6719), .ZN(n6805) );
NAND2_X1 U28768 ( .A1(n6785), .A2(n6786), .ZN(n14861) );
NOR2_X1 U28769 ( .A1(n6794), .A2(n6795), .ZN(n6785) );
NOR2_X1 U28770 ( .A1(n6787), .A2(n6788), .ZN(n6786) );
NOR2_X1 U28771 ( .A1(n10618), .A2(n6719), .ZN(n6795) );
NAND2_X1 U28772 ( .A1(n8136), .A2(n8137), .ZN(n15565) );
NOR2_X1 U28773 ( .A1(n8140), .A2(n7716), .ZN(n8136) );
NOR2_X1 U28774 ( .A1(n8138), .A2(n8139), .ZN(n8137) );
NOR2_X1 U28775 ( .A1(n11303), .A2(n20931), .ZN(n8140) );
NAND2_X1 U28776 ( .A1(n8131), .A2(n8132), .ZN(n15024) );
NOR2_X1 U28777 ( .A1(n8135), .A2(n7716), .ZN(n8131) );
NOR2_X1 U28778 ( .A1(n8133), .A2(n8134), .ZN(n8132) );
NOR2_X1 U28779 ( .A1(n10780), .A2(n16355), .ZN(n8135) );
NAND2_X1 U28780 ( .A1(n7895), .A2(n7896), .ZN(n15782) );
NOR2_X1 U28781 ( .A1(n7899), .A2(n7900), .ZN(n7895) );
NOR2_X1 U28782 ( .A1(n7897), .A2(n7898), .ZN(n7896) );
NOR2_X1 U28783 ( .A1(n11518), .A2(n16388), .ZN(n7900) );
NAND2_X1 U28784 ( .A1(n7913), .A2(n7914), .ZN(n15779) );
NOR2_X1 U28785 ( .A1(n7917), .A2(n7918), .ZN(n7913) );
NOR2_X1 U28786 ( .A1(n7915), .A2(n7916), .ZN(n7914) );
NOR2_X1 U28787 ( .A1(n11511), .A2(n16388), .ZN(n7918) );
NAND2_X1 U28788 ( .A1(n7919), .A2(n7920), .ZN(n15776) );
NOR2_X1 U28789 ( .A1(n7923), .A2(n7924), .ZN(n7919) );
NOR2_X1 U28790 ( .A1(n7921), .A2(n7922), .ZN(n7920) );
NOR2_X1 U28791 ( .A1(n11507), .A2(n16388), .ZN(n7924) );
NAND2_X1 U28792 ( .A1(n7979), .A2(n7980), .ZN(n15771) );
NOR2_X1 U28793 ( .A1(n7983), .A2(n7984), .ZN(n7979) );
NOR2_X1 U28794 ( .A1(n7981), .A2(n7982), .ZN(n7980) );
NOR2_X1 U28795 ( .A1(n11497), .A2(n7875), .ZN(n7984) );
NAND2_X1 U28796 ( .A1(n7991), .A2(n7992), .ZN(n15763) );
NOR2_X1 U28797 ( .A1(n7995), .A2(n7996), .ZN(n7991) );
NOR2_X1 U28798 ( .A1(n7993), .A2(n7994), .ZN(n7992) );
NOR2_X1 U28799 ( .A1(n11486), .A2(n7875), .ZN(n7996) );
NAND2_X1 U28800 ( .A1(n7943), .A2(n7944), .ZN(n15222) );
NOR2_X1 U28801 ( .A1(n7947), .A2(n7948), .ZN(n7943) );
NOR2_X1 U28802 ( .A1(n7945), .A2(n7946), .ZN(n7944) );
NOR2_X1 U28803 ( .A1(n10977), .A2(n7875), .ZN(n7948) );
NAND2_X1 U28804 ( .A1(n7949), .A2(n7950), .ZN(n15207) );
NOR2_X1 U28805 ( .A1(n7953), .A2(n7954), .ZN(n7949) );
NOR2_X1 U28806 ( .A1(n7951), .A2(n7952), .ZN(n7950) );
NOR2_X1 U28807 ( .A1(n10962), .A2(n7875), .ZN(n7954) );
NAND2_X1 U28808 ( .A1(n7955), .A2(n7956), .ZN(n15192) );
NOR2_X1 U28809 ( .A1(n7959), .A2(n7960), .ZN(n7955) );
NOR2_X1 U28810 ( .A1(n7957), .A2(n7958), .ZN(n7956) );
NOR2_X1 U28811 ( .A1(n10947), .A2(n7875), .ZN(n7960) );
NAND2_X1 U28812 ( .A1(n7961), .A2(n7962), .ZN(n15177) );
NOR2_X1 U28813 ( .A1(n7965), .A2(n7966), .ZN(n7961) );
NOR2_X1 U28814 ( .A1(n7963), .A2(n7964), .ZN(n7962) );
NOR2_X1 U28815 ( .A1(n10932), .A2(n7875), .ZN(n7966) );
NAND2_X1 U28816 ( .A1(n7967), .A2(n7968), .ZN(n15162) );
NOR2_X1 U28817 ( .A1(n7971), .A2(n7972), .ZN(n7967) );
NOR2_X1 U28818 ( .A1(n7969), .A2(n7970), .ZN(n7968) );
NOR2_X1 U28819 ( .A1(n10917), .A2(n7875), .ZN(n7972) );
NAND2_X1 U28820 ( .A1(n7973), .A2(n7974), .ZN(n15147) );
NOR2_X1 U28821 ( .A1(n7977), .A2(n7978), .ZN(n7973) );
NOR2_X1 U28822 ( .A1(n7975), .A2(n7976), .ZN(n7974) );
NOR2_X1 U28823 ( .A1(n10902), .A2(n7875), .ZN(n7978) );
NAND2_X1 U28824 ( .A1(n7985), .A2(n7986), .ZN(n15132) );
NOR2_X1 U28825 ( .A1(n7989), .A2(n7990), .ZN(n7985) );
NOR2_X1 U28826 ( .A1(n7987), .A2(n7988), .ZN(n7986) );
NOR2_X1 U28827 ( .A1(n10887), .A2(n7875), .ZN(n7990) );
NAND2_X1 U28828 ( .A1(n7997), .A2(n7998), .ZN(n15117) );
NOR2_X1 U28829 ( .A1(n8001), .A2(n8002), .ZN(n7997) );
NOR2_X1 U28830 ( .A1(n7999), .A2(n8000), .ZN(n7998) );
NOR2_X1 U28831 ( .A1(n10872), .A2(n7875), .ZN(n8002) );
NAND2_X1 U28832 ( .A1(n8003), .A2(n8004), .ZN(n15102) );
NOR2_X1 U28833 ( .A1(n8007), .A2(n8008), .ZN(n8003) );
NOR2_X1 U28834 ( .A1(n8005), .A2(n8006), .ZN(n8004) );
NOR2_X1 U28835 ( .A1(n10857), .A2(n7875), .ZN(n8008) );
NAND2_X1 U28836 ( .A1(n7867), .A2(n7868), .ZN(n14988) );
NOR2_X1 U28837 ( .A1(n7873), .A2(n7874), .ZN(n7867) );
NOR2_X1 U28838 ( .A1(n7869), .A2(n7870), .ZN(n7868) );
NOR2_X1 U28839 ( .A1(n10744), .A2(n16388), .ZN(n7874) );
NAND2_X1 U28840 ( .A1(n7877), .A2(n7878), .ZN(n14974) );
NOR2_X1 U28841 ( .A1(n7881), .A2(n7882), .ZN(n7877) );
NOR2_X1 U28842 ( .A1(n7879), .A2(n7880), .ZN(n7878) );
NOR2_X1 U28843 ( .A1(n10730), .A2(n16388), .ZN(n7882) );
NAND2_X1 U28844 ( .A1(n7889), .A2(n7890), .ZN(n14960) );
NOR2_X1 U28845 ( .A1(n7893), .A2(n7894), .ZN(n7889) );
NOR2_X1 U28846 ( .A1(n7891), .A2(n7892), .ZN(n7890) );
NOR2_X1 U28847 ( .A1(n10716), .A2(n16388), .ZN(n7894) );
NAND2_X1 U28848 ( .A1(n7901), .A2(n7902), .ZN(n14947) );
NOR2_X1 U28849 ( .A1(n7905), .A2(n7906), .ZN(n7901) );
NOR2_X1 U28850 ( .A1(n7903), .A2(n7904), .ZN(n7902) );
NOR2_X1 U28851 ( .A1(n10703), .A2(n16388), .ZN(n7906) );
NAND2_X1 U28852 ( .A1(n7883), .A2(n7884), .ZN(n14926) );
NOR2_X1 U28853 ( .A1(n7887), .A2(n7888), .ZN(n7883) );
NOR2_X1 U28854 ( .A1(n7885), .A2(n7886), .ZN(n7884) );
NOR2_X1 U28855 ( .A1(n10682), .A2(n16388), .ZN(n7888) );
NAND2_X1 U28856 ( .A1(n7907), .A2(n7908), .ZN(n14916) );
NOR2_X1 U28857 ( .A1(n7911), .A2(n7912), .ZN(n7907) );
NOR2_X1 U28858 ( .A1(n7909), .A2(n7910), .ZN(n7908) );
NOR2_X1 U28859 ( .A1(n10672), .A2(n16388), .ZN(n7912) );
NAND2_X1 U28860 ( .A1(n7925), .A2(n7926), .ZN(n14908) );
NOR2_X1 U28861 ( .A1(n7929), .A2(n7930), .ZN(n7925) );
NOR2_X1 U28862 ( .A1(n7927), .A2(n7928), .ZN(n7926) );
NOR2_X1 U28863 ( .A1(n10664), .A2(n16388), .ZN(n7930) );
NAND2_X1 U28864 ( .A1(n8009), .A2(n8010), .ZN(n14893) );
NOR2_X1 U28865 ( .A1(n8013), .A2(n8014), .ZN(n8009) );
NOR2_X1 U28866 ( .A1(n8011), .A2(n8012), .ZN(n8010) );
NOR2_X1 U28867 ( .A1(n10649), .A2(n7875), .ZN(n8014) );
NAND2_X1 U28868 ( .A1(n7937), .A2(n7938), .ZN(n14877) );
NOR2_X1 U28869 ( .A1(n7941), .A2(n7942), .ZN(n7937) );
NOR2_X1 U28870 ( .A1(n7939), .A2(n7940), .ZN(n7938) );
NOR2_X1 U28871 ( .A1(n10634), .A2(n16388), .ZN(n7942) );
NAND2_X1 U28872 ( .A1(n7931), .A2(n7932), .ZN(n14867) );
NOR2_X1 U28873 ( .A1(n7935), .A2(n7936), .ZN(n7931) );
NOR2_X1 U28874 ( .A1(n7933), .A2(n7934), .ZN(n7932) );
NOR2_X1 U28875 ( .A1(n10624), .A2(n16388), .ZN(n7936) );
NAND2_X1 U28876 ( .A1(n7061), .A2(n7062), .ZN(n15566) );
NOR2_X1 U28877 ( .A1(n7059), .A2(n7066), .ZN(n7061) );
NOR2_X1 U28878 ( .A1(n7063), .A2(n7064), .ZN(n7062) );
NOR2_X1 U28879 ( .A1(n11305), .A2(n7040), .ZN(n7066) );
NAND2_X1 U28880 ( .A1(n7053), .A2(n7054), .ZN(n15023) );
NOR2_X1 U28881 ( .A1(n7059), .A2(n7060), .ZN(n7053) );
NOR2_X1 U28882 ( .A1(n7055), .A2(n7056), .ZN(n7054) );
NOR2_X1 U28883 ( .A1(n10779), .A2(n7040), .ZN(n7060) );
NAND2_X1 U28884 ( .A1(n7372), .A2(n7373), .ZN(n15226) );
NOR2_X1 U28885 ( .A1(n7378), .A2(n7379), .ZN(n7372) );
NOR2_X1 U28886 ( .A1(n7374), .A2(n7375), .ZN(n7373) );
NOR2_X1 U28887 ( .A1(n10981), .A2(n16393), .ZN(n7379) );
NAND2_X1 U28888 ( .A1(n7548), .A2(n7549), .ZN(n15224) );
NOR2_X1 U28889 ( .A1(n7554), .A2(n7555), .ZN(n7548) );
NOR2_X1 U28890 ( .A1(n7550), .A2(n7551), .ZN(n7549) );
NOR2_X1 U28891 ( .A1(n11307), .A2(n7323), .ZN(n7554) );
NAND2_X1 U28892 ( .A1(n7412), .A2(n7413), .ZN(n15213) );
NOR2_X1 U28893 ( .A1(n7418), .A2(n7419), .ZN(n7412) );
NOR2_X1 U28894 ( .A1(n7414), .A2(n7415), .ZN(n7413) );
NOR2_X1 U28895 ( .A1(n10968), .A2(n16394), .ZN(n7419) );
NAND2_X1 U28896 ( .A1(n7420), .A2(n7421), .ZN(n15198) );
NOR2_X1 U28897 ( .A1(n7426), .A2(n7427), .ZN(n7420) );
NOR2_X1 U28898 ( .A1(n7422), .A2(n7423), .ZN(n7421) );
NOR2_X1 U28899 ( .A1(n10953), .A2(n16394), .ZN(n7427) );
NAND2_X1 U28900 ( .A1(n7428), .A2(n7429), .ZN(n15183) );
NOR2_X1 U28901 ( .A1(n7434), .A2(n7435), .ZN(n7428) );
NOR2_X1 U28902 ( .A1(n7430), .A2(n7431), .ZN(n7429) );
NOR2_X1 U28903 ( .A1(n10938), .A2(n16394), .ZN(n7435) );
NAND2_X1 U28904 ( .A1(n7436), .A2(n7437), .ZN(n15168) );
NOR2_X1 U28905 ( .A1(n7442), .A2(n7443), .ZN(n7436) );
NOR2_X1 U28906 ( .A1(n7438), .A2(n7439), .ZN(n7437) );
NOR2_X1 U28907 ( .A1(n10923), .A2(n16394), .ZN(n7443) );
NAND2_X1 U28908 ( .A1(n7444), .A2(n7445), .ZN(n15153) );
NOR2_X1 U28909 ( .A1(n7450), .A2(n7451), .ZN(n7444) );
NOR2_X1 U28910 ( .A1(n7446), .A2(n7447), .ZN(n7445) );
NOR2_X1 U28911 ( .A1(n10908), .A2(n16394), .ZN(n7451) );
NAND2_X1 U28912 ( .A1(n7452), .A2(n7453), .ZN(n15138) );
NOR2_X1 U28913 ( .A1(n7458), .A2(n7459), .ZN(n7452) );
NOR2_X1 U28914 ( .A1(n7454), .A2(n7455), .ZN(n7453) );
NOR2_X1 U28915 ( .A1(n10893), .A2(n16394), .ZN(n7459) );
NAND2_X1 U28916 ( .A1(n7468), .A2(n7469), .ZN(n15123) );
NOR2_X1 U28917 ( .A1(n7474), .A2(n7475), .ZN(n7468) );
NOR2_X1 U28918 ( .A1(n7470), .A2(n7471), .ZN(n7469) );
NOR2_X1 U28919 ( .A1(n10878), .A2(n16394), .ZN(n7475) );
NAND2_X1 U28920 ( .A1(n7484), .A2(n7485), .ZN(n15108) );
NOR2_X1 U28921 ( .A1(n7490), .A2(n7491), .ZN(n7484) );
NOR2_X1 U28922 ( .A1(n7486), .A2(n7487), .ZN(n7485) );
NOR2_X1 U28923 ( .A1(n10863), .A2(n16394), .ZN(n7491) );
NAND2_X1 U28924 ( .A1(n7492), .A2(n7493), .ZN(n15091) );
NOR2_X1 U28925 ( .A1(n7498), .A2(n7499), .ZN(n7492) );
NOR2_X1 U28926 ( .A1(n7494), .A2(n7495), .ZN(n7493) );
NOR2_X1 U28927 ( .A1(n10846), .A2(n16394), .ZN(n7499) );
NAND2_X1 U28928 ( .A1(n7508), .A2(n7509), .ZN(n15076) );
NOR2_X1 U28929 ( .A1(n7514), .A2(n7515), .ZN(n7508) );
NOR2_X1 U28930 ( .A1(n7510), .A2(n7511), .ZN(n7509) );
NOR2_X1 U28931 ( .A1(n10832), .A2(n16392), .ZN(n7514) );
NAND2_X1 U28932 ( .A1(n7516), .A2(n7517), .ZN(n15061) );
NOR2_X1 U28933 ( .A1(n7522), .A2(n7523), .ZN(n7516) );
NOR2_X1 U28934 ( .A1(n7518), .A2(n7519), .ZN(n7517) );
NOR2_X1 U28935 ( .A1(n10817), .A2(n7323), .ZN(n7522) );
NAND2_X1 U28936 ( .A1(n7524), .A2(n7525), .ZN(n15047) );
NOR2_X1 U28937 ( .A1(n7530), .A2(n7531), .ZN(n7524) );
NOR2_X1 U28938 ( .A1(n7526), .A2(n7527), .ZN(n7525) );
NOR2_X1 U28939 ( .A1(n10803), .A2(n16392), .ZN(n7530) );
NAND2_X1 U28940 ( .A1(n7532), .A2(n7533), .ZN(n15032) );
NOR2_X1 U28941 ( .A1(n7538), .A2(n7539), .ZN(n7532) );
NOR2_X1 U28942 ( .A1(n7534), .A2(n7535), .ZN(n7533) );
NOR2_X1 U28943 ( .A1(n10788), .A2(n7323), .ZN(n7538) );
NAND2_X1 U28944 ( .A1(n7540), .A2(n7541), .ZN(n15011) );
NOR2_X1 U28945 ( .A1(n7546), .A2(n7547), .ZN(n7540) );
NOR2_X1 U28946 ( .A1(n7542), .A2(n7543), .ZN(n7541) );
NOR2_X1 U28947 ( .A1(n10769), .A2(n16392), .ZN(n7546) );
NAND2_X1 U28948 ( .A1(n7556), .A2(n7557), .ZN(n14997) );
NOR2_X1 U28949 ( .A1(n7565), .A2(n7566), .ZN(n7556) );
NOR2_X1 U28950 ( .A1(n7558), .A2(n7559), .ZN(n7557) );
NOR2_X1 U28951 ( .A1(n10759), .A2(n7323), .ZN(n7565) );
NAND2_X1 U28952 ( .A1(n7324), .A2(n7325), .ZN(n14969) );
NOR2_X1 U28953 ( .A1(n7330), .A2(n7331), .ZN(n7324) );
NOR2_X1 U28954 ( .A1(n7326), .A2(n7327), .ZN(n7325) );
NOR2_X1 U28955 ( .A1(n10725), .A2(n16393), .ZN(n7331) );
NAND2_X1 U28956 ( .A1(n7340), .A2(n7341), .ZN(n14955) );
NOR2_X1 U28957 ( .A1(n7346), .A2(n7347), .ZN(n7340) );
NOR2_X1 U28958 ( .A1(n7342), .A2(n7343), .ZN(n7341) );
NOR2_X1 U28959 ( .A1(n10711), .A2(n16393), .ZN(n7347) );
NAND2_X1 U28960 ( .A1(n7356), .A2(n7357), .ZN(n14942) );
NOR2_X1 U28961 ( .A1(n7362), .A2(n7363), .ZN(n7356) );
NOR2_X1 U28962 ( .A1(n7358), .A2(n7359), .ZN(n7357) );
NOR2_X1 U28963 ( .A1(n10698), .A2(n16393), .ZN(n7363) );
NAND2_X1 U28964 ( .A1(n7332), .A2(n7333), .ZN(n14923) );
NOR2_X1 U28965 ( .A1(n7338), .A2(n7339), .ZN(n7332) );
NOR2_X1 U28966 ( .A1(n7334), .A2(n7335), .ZN(n7333) );
NOR2_X1 U28967 ( .A1(n10679), .A2(n16393), .ZN(n7339) );
NAND2_X1 U28968 ( .A1(n7364), .A2(n7365), .ZN(n14913) );
NOR2_X1 U28969 ( .A1(n7370), .A2(n7371), .ZN(n7364) );
NOR2_X1 U28970 ( .A1(n7366), .A2(n7367), .ZN(n7365) );
NOR2_X1 U28971 ( .A1(n10669), .A2(n16393), .ZN(n7371) );
NAND2_X1 U28972 ( .A1(n7388), .A2(n7389), .ZN(n14905) );
NOR2_X1 U28973 ( .A1(n7394), .A2(n7395), .ZN(n7388) );
NOR2_X1 U28974 ( .A1(n7390), .A2(n7391), .ZN(n7389) );
NOR2_X1 U28975 ( .A1(n10661), .A2(n16393), .ZN(n7395) );
NAND2_X1 U28976 ( .A1(n7500), .A2(n7501), .ZN(n14890) );
NOR2_X1 U28977 ( .A1(n7506), .A2(n7507), .ZN(n7500) );
NOR2_X1 U28978 ( .A1(n7502), .A2(n7503), .ZN(n7501) );
NOR2_X1 U28979 ( .A1(n10646), .A2(n16394), .ZN(n7507) );
NAND2_X1 U28980 ( .A1(n7476), .A2(n7477), .ZN(n14887) );
NOR2_X1 U28981 ( .A1(n7482), .A2(n7483), .ZN(n7476) );
NOR2_X1 U28982 ( .A1(n7478), .A2(n7479), .ZN(n7477) );
NOR2_X1 U28983 ( .A1(n10644), .A2(n16394), .ZN(n7483) );
NAND2_X1 U28984 ( .A1(n7404), .A2(n7405), .ZN(n14874) );
NOR2_X1 U28985 ( .A1(n7410), .A2(n7411), .ZN(n7404) );
NOR2_X1 U28986 ( .A1(n7406), .A2(n7407), .ZN(n7405) );
NOR2_X1 U28987 ( .A1(n10631), .A2(n16393), .ZN(n7411) );
NAND2_X1 U28988 ( .A1(n7396), .A2(n7397), .ZN(n14864) );
NOR2_X1 U28989 ( .A1(n7402), .A2(n7403), .ZN(n7396) );
NOR2_X1 U28990 ( .A1(n7398), .A2(n7399), .ZN(n7397) );
NOR2_X1 U28991 ( .A1(n10621), .A2(n16393), .ZN(n7403) );
NAND2_X1 U28992 ( .A1(n7460), .A2(n7461), .ZN(n14860) );
NOR2_X1 U28993 ( .A1(n7466), .A2(n7467), .ZN(n7460) );
NOR2_X1 U28994 ( .A1(n7462), .A2(n7463), .ZN(n7461) );
NOR2_X1 U28995 ( .A1(n10617), .A2(n16394), .ZN(n7467) );
NAND2_X1 U28996 ( .A1(n7380), .A2(n7381), .ZN(n14858) );
NOR2_X1 U28997 ( .A1(n7386), .A2(n7387), .ZN(n7380) );
NOR2_X1 U28998 ( .A1(n7382), .A2(n7383), .ZN(n7381) );
NOR2_X1 U28999 ( .A1(n10615), .A2(n16393), .ZN(n7387) );
NAND2_X1 U29000 ( .A1(n7348), .A2(n7349), .ZN(n14853) );
NOR2_X1 U29001 ( .A1(n7354), .A2(n7355), .ZN(n7348) );
NOR2_X1 U29002 ( .A1(n7350), .A2(n7351), .ZN(n7349) );
NOR2_X1 U29003 ( .A1(n10610), .A2(n16393), .ZN(n7355) );
NAND2_X1 U29004 ( .A1(n7312), .A2(n7313), .ZN(n14983) );
NOR2_X1 U29005 ( .A1(n7320), .A2(n7321), .ZN(n7312) );
NOR2_X1 U29006 ( .A1(n7314), .A2(n7315), .ZN(n7313) );
NOR2_X1 U29007 ( .A1(n10739), .A2(n16393), .ZN(n7321) );
NAND2_X1 U29008 ( .A1(n2096), .A2(n2097), .ZN(n15577) );
NOR2_X1 U29009 ( .A1(n2114), .A2(n2115), .ZN(n2096) );
NOR2_X1 U29010 ( .A1(n2098), .A2(n2099), .ZN(n2097) );
NOR2_X1 U29011 ( .A1(n11311), .A2(n16453), .ZN(n2115) );
NAND2_X1 U29012 ( .A1(n2173), .A2(n2174), .ZN(n15595) );
NOR2_X1 U29013 ( .A1(n2185), .A2(n2186), .ZN(n2173) );
NOR2_X1 U29014 ( .A1(n2175), .A2(n2176), .ZN(n2174) );
NOR2_X1 U29015 ( .A1(n11323), .A2(n16450), .ZN(n2186) );
NAND2_X1 U29016 ( .A1(n7042), .A2(n7043), .ZN(n15572) );
NOR2_X1 U29017 ( .A1(n7050), .A2(n7051), .ZN(n7042) );
NOR2_X1 U29018 ( .A1(n7044), .A2(n7045), .ZN(n7043) );
NOR2_X1 U29019 ( .A1(n11476), .A2(n7040), .ZN(n7051) );
NAND2_X1 U29020 ( .A1(n7015), .A2(n7016), .ZN(n15255) );
AND2_X1 U29021 ( .A1(n7017), .A2(n7018), .ZN(n7016) );
NOR2_X1 U29022 ( .A1(n7026), .A2(n7027), .ZN(n7015) );
NAND2_X1 U29023 ( .A1(crash_dump_o_96_), .A2(n16403), .ZN(n7018) );
INV_X1 U29024 ( .A(n22961), .ZN(n16328) );
INV_X1 U29025 ( .A(n24098), .ZN(n20163) );
INV_X1 U29026 ( .A(n23651), .ZN(n20312) );
INV_X1 U29027 ( .A(n23378), .ZN(n20465) );
INV_X1 U29028 ( .A(n23512), .ZN(n20388) );
INV_X1 U29029 ( .A(n23954), .ZN(n20079) );
INV_X1 U29030 ( .A(n22670), .ZN(n20662) );
INV_X1 U29031 ( .A(n22793), .ZN(n16329) );
INV_X1 U29032 ( .A(n22776), .ZN(n20628) );
INV_X1 U29033 ( .A(n23939), .ZN(n16330) );
INV_X1 U29034 ( .A(n23939), .ZN(n20165) );
INV_X1 U29035 ( .A(n22944), .ZN(n20624) );
BUF_X1 U29036 ( .A(n20241), .Z(n16331) );
BUF_X1 U29037 ( .A(n20392), .Z(n16332) );
BUF_X1 U29038 ( .A(n20473), .Z(n16333) );
INV_X1 U29039 ( .A(n23480), .ZN(n20241) );
INV_X1 U29040 ( .A(n23223), .ZN(n20392) );
INV_X1 U29041 ( .A(n23112), .ZN(n20473) );
NAND2_X1 U29042 ( .A1(n352), .A2(n353), .ZN(rf_wdata_wb_ecc_o_31_) );
NOR2_X1 U29043 ( .A1(n379), .A2(n380), .ZN(n352) );
NAND2_X1 U29044 ( .A1(n388), .A2(n389), .ZN(n379) );
NOR2_X1 U29045 ( .A1(n390), .A2(n391), .ZN(n389) );
AND2_X1 U29046 ( .A1(n20820), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_31), .ZN(n390) );
NAND2_X1 U29047 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
NAND2_X1 U29048 ( .A1(n1409), .A2(n1410), .ZN(n1408) );
NAND2_X1 U29049 ( .A1(ex_block_i_alu_i_adder_in_b_29), .A2(n21233), .ZN(n21234) );
NAND2_X1 U29050 ( .A1(ex_block_i_alu_i_adder_in_b_30), .A2(n21242), .ZN(n21243) );
NAND2_X1 U29051 ( .A1(ex_block_i_alu_i_adder_in_b_25), .A2(n21191), .ZN(n21192) );
NAND2_X1 U29052 ( .A1(ex_block_i_alu_i_adder_in_b_26), .A2(n21200), .ZN(n21201) );
NAND2_X1 U29053 ( .A1(ex_block_i_alu_i_adder_in_b_22), .A2(n21164), .ZN(n21165) );
NAND2_X1 U29054 ( .A1(ex_block_i_alu_i_adder_in_b_23), .A2(n21173), .ZN(n21174) );
NAND2_X1 U29055 ( .A1(ex_block_i_alu_i_adder_in_b_19), .A2(n21137), .ZN(n21138) );
NAND2_X1 U29056 ( .A1(ex_block_i_alu_i_adder_in_b_20), .A2(n21146), .ZN(n21147) );
NAND2_X1 U29057 ( .A1(ex_block_i_alu_i_adder_in_b_15), .A2(n21096), .ZN(n21097) );
NAND2_X1 U29058 ( .A1(ex_block_i_alu_i_adder_in_b_16), .A2(n21105), .ZN(n21106) );
NAND2_X1 U29059 ( .A1(ex_block_i_alu_i_adder_in_b_12), .A2(n21069), .ZN(n21070) );
NAND2_X1 U29060 ( .A1(ex_block_i_alu_i_adder_in_b_13), .A2(n21078), .ZN(n21079) );
NAND2_X1 U29061 ( .A1(ex_block_i_alu_i_adder_in_b_9), .A2(n21042), .ZN(n21043) );
NAND2_X1 U29062 ( .A1(ex_block_i_alu_i_adder_in_b_10), .A2(n21051), .ZN(n21052) );
NAND2_X1 U29063 ( .A1(ex_block_i_alu_i_adder_in_b_5), .A2(n21030), .ZN(n21031) );
NAND2_X1 U29064 ( .A1(ex_block_i_alu_i_adder_in_b_6), .A2(n21033), .ZN(n21034) );
NAND2_X1 U29065 ( .A1(ex_block_i_alu_i_adder_in_b_2), .A2(n21021), .ZN(n21022) );
NAND2_X1 U29066 ( .A1(ex_block_i_alu_i_adder_in_b_3), .A2(n21024), .ZN(n21025) );
NOR2_X1 U29067 ( .A1(n16364), .A2(n20760), .ZN(n9961) );
NAND2_X1 U29068 ( .A1(n21632), .A2(n21631), .ZN(n21648) );
NOR2_X1 U29069 ( .A1(n9961), .A2(n9962), .ZN(n9960) );
NOR2_X1 U29070 ( .A1(n21256), .A2(n21257), .ZN(n21259) );
BUF_X1 U29071 ( .A(n16336), .Z(n16337) );
BUF_X1 U29072 ( .A(n16336), .Z(n16338) );
BUF_X1 U29073 ( .A(n16336), .Z(n16339) );
BUF_X1 U29074 ( .A(n16336), .Z(n16340) );
BUF_X1 U29075 ( .A(n16336), .Z(n16341) );
BUF_X1 U29076 ( .A(n16336), .Z(n16342) );
BUF_X1 U29077 ( .A(n16336), .Z(n16343) );
BUF_X1 U29078 ( .A(n19748), .Z(n16344) );
BUF_X1 U29079 ( .A(n20924), .Z(n16354) );
BUF_X1 U29080 ( .A(n22014), .Z(n16359) );
BUF_X1 U29081 ( .A(n22015), .Z(n16360) );
INV_X1 U29082 ( .A(n16366), .ZN(n16365) );
INV_X1 U29083 ( .A(n16386), .ZN(n16385) );
BUF_X1 U29084 ( .A(n4275), .Z(n16423) );
BUF_X1 U29085 ( .A(n3061), .Z(n16437) );
BUF_X1 U29086 ( .A(n3061), .Z(n16438) );
BUF_X1 U29087 ( .A(n2901), .Z(n16443) );
BUF_X1 U29088 ( .A(n2900), .Z(n16444) );
INV_X1 U29089 ( .A(n16447), .ZN(n16446) );
INV_X1 U29090 ( .A(n16449), .ZN(n16448) );
INV_X1 U29091 ( .A(n16467), .ZN(n16466) );
INV_X4 U32362 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_sign_a), .ZN(n20084) );
INV_X4 U32363 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_sign_b), .ZN(n20762) );
NOR2_X4 U32364 ( .A1(n16200), .A2(n20804), .ZN(n22546) );
NOR2_X4 U32365 ( .A1(n20807), .A2(n20675), .ZN(n25258) );
NAND2_X4 U32366 ( .A1(n22546), .A2(n25258), .ZN(n23046) );
NAND2_X4 U32367 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n22547) );
NAND2_X4 U32368 ( .A1(n20674), .A2(n22547), .ZN(n22549) );
NAND2_X4 U32369 ( .A1(n20640), .A2(n23046), .ZN(n22548) );
NAND2_X4 U32370 ( .A1(n22549), .A2(n22548), .ZN(n22553) );
NAND2_X4 U32371 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n22550) );
NOR2_X4 U32372 ( .A1(n20804), .A2(n20675), .ZN(n22875) );
OR2_X4 U32373 ( .A1(n22550), .A2(n22875), .ZN(n22552) );
NAND2_X4 U32374 ( .A1(n22875), .A2(n22550), .ZN(n22551) );
NAND2_X4 U32375 ( .A1(n22552), .A2(n22551), .ZN(n23045) );
NAND2_X4 U32376 ( .A1(n22553), .A2(n20671), .ZN(n22555) );
OR2_X4 U32377 ( .A1(n20671), .A2(n22553), .ZN(n22554) );
NAND2_X4 U32378 ( .A1(n22555), .A2(n22554), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N37) );
NAND2_X4 U32379 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n22821) );
NAND2_X4 U32380 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n22692) );
NAND2_X4 U32381 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n22607) );
NAND2_X4 U32382 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n22567) );
NAND2_X4 U32383 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n22583) );
NOR2_X4 U32384 ( .A1(n16200), .A2(n20789), .ZN(n22556) );
NOR2_X4 U32385 ( .A1(n20792), .A2(n20675), .ZN(n22569) );
NAND2_X4 U32386 ( .A1(n22556), .A2(n22569), .ZN(n22557) );
NAND2_X4 U32387 ( .A1(n20637), .A2(n22557), .ZN(n22559) );
NAND2_X4 U32388 ( .A1(n20669), .A2(n22583), .ZN(n22558) );
NAND2_X4 U32389 ( .A1(n22559), .A2(n22558), .ZN(n22563) );
NAND2_X4 U32390 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n22560) );
NOR2_X4 U32391 ( .A1(n20789), .A2(n20675), .ZN(n22589) );
OR2_X4 U32392 ( .A1(n22560), .A2(n22589), .ZN(n22562) );
NAND2_X4 U32393 ( .A1(n22589), .A2(n22560), .ZN(n22561) );
NAND2_X4 U32394 ( .A1(n22562), .A2(n22561), .ZN(n22582) );
NAND2_X4 U32395 ( .A1(n22563), .A2(n20667), .ZN(n22565) );
OR2_X4 U32396 ( .A1(n20667), .A2(n22563), .ZN(n22564) );
NAND2_X4 U32397 ( .A1(n22565), .A2(n22564), .ZN(n22566) );
NAND2_X4 U32398 ( .A1(n20602), .A2(n22566), .ZN(n22579) );
NAND2_X4 U32399 ( .A1(n20636), .A2(n22567), .ZN(n22577) );
NAND2_X4 U32400 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n22617) );
NAND2_X4 U32401 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n22568) );
OR2_X4 U32402 ( .A1(n22568), .A2(n22569), .ZN(n22571) );
NAND2_X4 U32403 ( .A1(n22569), .A2(n22568), .ZN(n22570) );
NAND2_X4 U32404 ( .A1(n22571), .A2(n22570), .ZN(n22573) );
NAND2_X4 U32405 ( .A1(n20635), .A2(n22573), .ZN(n22576) );
NOR2_X4 U32406 ( .A1(n16200), .A2(n20792), .ZN(n22572) );
NOR2_X4 U32407 ( .A1(n20795), .A2(n20675), .ZN(n22626) );
NAND2_X4 U32408 ( .A1(n22572), .A2(n22626), .ZN(n22616) );
NAND2_X4 U32409 ( .A1(n20668), .A2(n22617), .ZN(n22574) );
NAND2_X4 U32410 ( .A1(n20665), .A2(n22574), .ZN(n22575) );
NAND2_X4 U32411 ( .A1(n22576), .A2(n22575), .ZN(n22608) );
NAND2_X4 U32412 ( .A1(n22577), .A2(n22608), .ZN(n22578) );
NAND2_X4 U32413 ( .A1(n22579), .A2(n22578), .ZN(n22647) );
NAND2_X4 U32414 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n22645) );
OR2_X4 U32415 ( .A1(n22647), .A2(n20562), .ZN(n22581) );
NAND2_X4 U32416 ( .A1(n20562), .A2(n22647), .ZN(n22580) );
NAND2_X4 U32417 ( .A1(n22581), .A2(n22580), .ZN(n22603) );
NAND2_X4 U32418 ( .A1(n20637), .A2(n22582), .ZN(n22586) );
NAND2_X4 U32419 ( .A1(n20667), .A2(n22583), .ZN(n22584) );
NAND2_X4 U32420 ( .A1(n20669), .A2(n22584), .ZN(n22585) );
NAND2_X4 U32421 ( .A1(n22586), .A2(n22585), .ZN(n22655) );
NAND2_X4 U32422 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n22654) );
OR2_X4 U32423 ( .A1(n22655), .A2(n20600), .ZN(n22588) );
NAND2_X4 U32424 ( .A1(n20600), .A2(n22655), .ZN(n22587) );
NAND2_X4 U32425 ( .A1(n22588), .A2(n22587), .ZN(n22600) );
NAND2_X4 U32426 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n22662) );
NOR2_X4 U32427 ( .A1(n16200), .A2(n20786), .ZN(n22590) );
NAND2_X4 U32428 ( .A1(n22590), .A2(n22589), .ZN(n22591) );
NAND2_X4 U32429 ( .A1(n20633), .A2(n22591), .ZN(n22593) );
NAND2_X4 U32430 ( .A1(n20666), .A2(n22662), .ZN(n22592) );
NAND2_X4 U32431 ( .A1(n22593), .A2(n22592), .ZN(n22597) );
NAND2_X4 U32432 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n22594) );
NOR2_X4 U32433 ( .A1(n20786), .A2(n20675), .ZN(n22668) );
OR2_X4 U32434 ( .A1(n22594), .A2(n22668), .ZN(n22596) );
NAND2_X4 U32435 ( .A1(n22668), .A2(n22594), .ZN(n22595) );
NAND2_X4 U32436 ( .A1(n22596), .A2(n22595), .ZN(n22661) );
NAND2_X4 U32437 ( .A1(n22597), .A2(n20663), .ZN(n22599) );
OR2_X4 U32438 ( .A1(n20663), .A2(n22597), .ZN(n22598) );
NAND2_X4 U32439 ( .A1(n22599), .A2(n22598), .ZN(n22653) );
NAND2_X4 U32440 ( .A1(n22600), .A2(n20632), .ZN(n22602) );
OR2_X4 U32441 ( .A1(n20632), .A2(n22600), .ZN(n22601) );
NAND2_X4 U32442 ( .A1(n22602), .A2(n22601), .ZN(n22646) );
NAND2_X4 U32443 ( .A1(n22603), .A2(n20599), .ZN(n22605) );
OR2_X4 U32444 ( .A1(n20599), .A2(n22603), .ZN(n22604) );
NAND2_X4 U32445 ( .A1(n22605), .A2(n22604), .ZN(n22606) );
NAND2_X4 U32446 ( .A1(n20522), .A2(n22606), .ZN(n22642) );
NAND2_X4 U32447 ( .A1(n20561), .A2(n22607), .ZN(n22640) );
NAND2_X4 U32448 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n22614) );
OR2_X4 U32449 ( .A1(n22608), .A2(n20602), .ZN(n22610) );
NAND2_X4 U32450 ( .A1(n20602), .A2(n22608), .ZN(n22609) );
NAND2_X4 U32451 ( .A1(n22610), .A2(n22609), .ZN(n22611) );
NAND2_X4 U32452 ( .A1(n22611), .A2(n20636), .ZN(n22613) );
OR2_X4 U32453 ( .A1(n20636), .A2(n22611), .ZN(n22612) );
NAND2_X4 U32454 ( .A1(n22613), .A2(n22612), .ZN(n22615) );
NAND2_X4 U32455 ( .A1(n20560), .A2(n20601), .ZN(n22639) );
NAND2_X4 U32456 ( .A1(n22615), .A2(n22614), .ZN(n22637) );
NAND2_X4 U32457 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n22624) );
NAND2_X4 U32458 ( .A1(n20635), .A2(n22616), .ZN(n22619) );
NAND2_X4 U32459 ( .A1(n20665), .A2(n22617), .ZN(n22618) );
NAND2_X4 U32460 ( .A1(n22619), .A2(n22618), .ZN(n22620) );
NAND2_X4 U32461 ( .A1(n22620), .A2(n20668), .ZN(n22622) );
OR2_X4 U32462 ( .A1(n20668), .A2(n22620), .ZN(n22621) );
NAND2_X4 U32463 ( .A1(n22622), .A2(n22621), .ZN(n22623) );
NAND2_X4 U32464 ( .A1(n20598), .A2(n22623), .ZN(n22636) );
NAND2_X4 U32465 ( .A1(n20634), .A2(n22624), .ZN(n22634) );
NAND2_X4 U32466 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n22718) );
NAND2_X4 U32467 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n22625) );
OR2_X4 U32468 ( .A1(n22625), .A2(n22626), .ZN(n22628) );
NAND2_X4 U32469 ( .A1(n22626), .A2(n22625), .ZN(n22627) );
NAND2_X4 U32470 ( .A1(n22628), .A2(n22627), .ZN(n22630) );
NAND2_X4 U32471 ( .A1(n20631), .A2(n22630), .ZN(n22633) );
NOR2_X4 U32472 ( .A1(n16200), .A2(n20795), .ZN(n22629) );
NOR2_X4 U32473 ( .A1(n20798), .A2(n20675), .ZN(n22727) );
NAND2_X4 U32474 ( .A1(n22629), .A2(n22727), .ZN(n22717) );
NAND2_X4 U32475 ( .A1(n20664), .A2(n22718), .ZN(n22631) );
NAND2_X4 U32476 ( .A1(n20661), .A2(n22631), .ZN(n22632) );
NAND2_X4 U32477 ( .A1(n22633), .A2(n22632), .ZN(n22709) );
NAND2_X4 U32478 ( .A1(n22634), .A2(n22709), .ZN(n22635) );
NAND2_X4 U32479 ( .A1(n22636), .A2(n22635), .ZN(n22701) );
NAND2_X4 U32480 ( .A1(n22637), .A2(n22701), .ZN(n22638) );
NAND2_X4 U32481 ( .A1(n22639), .A2(n22638), .ZN(n22693) );
NAND2_X4 U32482 ( .A1(n22640), .A2(n22693), .ZN(n22641) );
NAND2_X4 U32483 ( .A1(n22642), .A2(n22641), .ZN(n22754) );
NAND2_X4 U32484 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n22752) );
OR2_X4 U32485 ( .A1(n22754), .A2(n20482), .ZN(n22644) );
NAND2_X4 U32486 ( .A1(n20482), .A2(n22754), .ZN(n22643) );
NAND2_X4 U32487 ( .A1(n22644), .A2(n22643), .ZN(n22688) );
NAND2_X4 U32488 ( .A1(n20562), .A2(n20599), .ZN(n22650) );
NAND2_X4 U32489 ( .A1(n22646), .A2(n22645), .ZN(n22648) );
NAND2_X4 U32490 ( .A1(n22648), .A2(n22647), .ZN(n22649) );
NAND2_X4 U32491 ( .A1(n22650), .A2(n22649), .ZN(n22762) );
NAND2_X4 U32492 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n22761) );
OR2_X4 U32493 ( .A1(n22762), .A2(n20520), .ZN(n22652) );
NAND2_X4 U32494 ( .A1(n20520), .A2(n22762), .ZN(n22651) );
NAND2_X4 U32495 ( .A1(n22652), .A2(n22651), .ZN(n22685) );
NAND2_X4 U32496 ( .A1(n20600), .A2(n22653), .ZN(n22658) );
NAND2_X4 U32497 ( .A1(n20632), .A2(n22654), .ZN(n22656) );
NAND2_X4 U32498 ( .A1(n22656), .A2(n22655), .ZN(n22657) );
NAND2_X4 U32499 ( .A1(n22658), .A2(n22657), .ZN(n22770) );
NAND2_X4 U32500 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n22768) );
OR2_X4 U32501 ( .A1(n22770), .A2(n20558), .ZN(n22660) );
NAND2_X4 U32502 ( .A1(n20558), .A2(n22770), .ZN(n22659) );
NAND2_X4 U32503 ( .A1(n22660), .A2(n22659), .ZN(n22682) );
NAND2_X4 U32504 ( .A1(n20633), .A2(n22661), .ZN(n22665) );
NAND2_X4 U32505 ( .A1(n20663), .A2(n22662), .ZN(n22663) );
NAND2_X4 U32506 ( .A1(n20666), .A2(n22663), .ZN(n22664) );
NAND2_X4 U32507 ( .A1(n22665), .A2(n22664), .ZN(n22778) );
NAND2_X4 U32508 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n22777) );
OR2_X4 U32509 ( .A1(n22778), .A2(n20596), .ZN(n22667) );
NAND2_X4 U32510 ( .A1(n20596), .A2(n22778), .ZN(n22666) );
NAND2_X4 U32511 ( .A1(n22667), .A2(n22666), .ZN(n22679) );
NAND2_X4 U32512 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n22785) );
NOR2_X4 U32513 ( .A1(n20683), .A2(n20783), .ZN(n22669) );
NAND2_X4 U32514 ( .A1(n22669), .A2(n22668), .ZN(n22670) );
NAND2_X4 U32515 ( .A1(n20629), .A2(n22670), .ZN(n22672) );
NAND2_X4 U32516 ( .A1(n20662), .A2(n22785), .ZN(n22671) );
NAND2_X4 U32517 ( .A1(n22672), .A2(n22671), .ZN(n22676) );
NAND2_X4 U32518 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n22673) );
NOR2_X4 U32519 ( .A1(n20783), .A2(n20675), .ZN(n22791) );
OR2_X4 U32520 ( .A1(n22673), .A2(n22791), .ZN(n22675) );
NAND2_X4 U32521 ( .A1(n22791), .A2(n22673), .ZN(n22674) );
NAND2_X4 U32522 ( .A1(n22675), .A2(n22674), .ZN(n22784) );
NAND2_X4 U32523 ( .A1(n22676), .A2(n20659), .ZN(n22678) );
OR2_X4 U32524 ( .A1(n20659), .A2(n22676), .ZN(n22677) );
NAND2_X4 U32525 ( .A1(n22678), .A2(n22677), .ZN(n22776) );
NAND2_X4 U32526 ( .A1(n22679), .A2(n20628), .ZN(n22681) );
OR2_X4 U32527 ( .A1(n20628), .A2(n22679), .ZN(n22680) );
NAND2_X4 U32528 ( .A1(n22681), .A2(n22680), .ZN(n22769) );
NAND2_X4 U32529 ( .A1(n22682), .A2(n20595), .ZN(n22684) );
OR2_X4 U32530 ( .A1(n20595), .A2(n22682), .ZN(n22683) );
NAND2_X4 U32531 ( .A1(n22684), .A2(n22683), .ZN(n22760) );
NAND2_X4 U32532 ( .A1(n22685), .A2(n20557), .ZN(n22687) );
OR2_X4 U32533 ( .A1(n20557), .A2(n22685), .ZN(n22686) );
NAND2_X4 U32534 ( .A1(n22687), .A2(n22686), .ZN(n22753) );
NAND2_X4 U32535 ( .A1(n22688), .A2(n20519), .ZN(n22690) );
OR2_X4 U32536 ( .A1(n20519), .A2(n22688), .ZN(n22689) );
NAND2_X4 U32537 ( .A1(n22690), .A2(n22689), .ZN(n22691) );
NAND2_X4 U32538 ( .A1(n20442), .A2(n22691), .ZN(n22749) );
NAND2_X4 U32539 ( .A1(n20481), .A2(n22692), .ZN(n22747) );
NAND2_X4 U32540 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n22699) );
OR2_X4 U32541 ( .A1(n22693), .A2(n20522), .ZN(n22695) );
NAND2_X4 U32542 ( .A1(n20522), .A2(n22693), .ZN(n22694) );
NAND2_X4 U32543 ( .A1(n22695), .A2(n22694), .ZN(n22696) );
NAND2_X4 U32544 ( .A1(n22696), .A2(n20561), .ZN(n22698) );
OR2_X4 U32545 ( .A1(n20561), .A2(n22696), .ZN(n22697) );
NAND2_X4 U32546 ( .A1(n22698), .A2(n22697), .ZN(n22700) );
NAND2_X4 U32547 ( .A1(n20480), .A2(n20521), .ZN(n22746) );
NAND2_X4 U32548 ( .A1(n22700), .A2(n22699), .ZN(n22744) );
NAND2_X4 U32549 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n22708) );
OR2_X4 U32550 ( .A1(n22701), .A2(n20560), .ZN(n22703) );
NAND2_X4 U32551 ( .A1(n20560), .A2(n22701), .ZN(n22702) );
NAND2_X4 U32552 ( .A1(n22703), .A2(n22702), .ZN(n22704) );
NAND2_X4 U32553 ( .A1(n22704), .A2(n20601), .ZN(n22706) );
OR2_X4 U32554 ( .A1(n20601), .A2(n22704), .ZN(n22705) );
NAND2_X4 U32555 ( .A1(n22706), .A2(n22705), .ZN(n22707) );
NAND2_X4 U32556 ( .A1(n20518), .A2(n22707), .ZN(n22743) );
NAND2_X4 U32557 ( .A1(n20559), .A2(n22708), .ZN(n22741) );
NAND2_X4 U32558 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n22715) );
OR2_X4 U32559 ( .A1(n22709), .A2(n20598), .ZN(n22711) );
NAND2_X4 U32560 ( .A1(n20598), .A2(n22709), .ZN(n22710) );
NAND2_X4 U32561 ( .A1(n22711), .A2(n22710), .ZN(n22712) );
NAND2_X4 U32562 ( .A1(n22712), .A2(n20634), .ZN(n22714) );
OR2_X4 U32563 ( .A1(n20634), .A2(n22712), .ZN(n22713) );
NAND2_X4 U32564 ( .A1(n22714), .A2(n22713), .ZN(n22716) );
NAND2_X4 U32565 ( .A1(n20556), .A2(n20597), .ZN(n22740) );
NAND2_X4 U32566 ( .A1(n22716), .A2(n22715), .ZN(n22738) );
NAND2_X4 U32567 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n22725) );
NAND2_X4 U32568 ( .A1(n20631), .A2(n22717), .ZN(n22720) );
NAND2_X4 U32569 ( .A1(n20661), .A2(n22718), .ZN(n22719) );
NAND2_X4 U32570 ( .A1(n22720), .A2(n22719), .ZN(n22721) );
NAND2_X4 U32571 ( .A1(n22721), .A2(n20664), .ZN(n22723) );
OR2_X4 U32572 ( .A1(n20664), .A2(n22721), .ZN(n22722) );
NAND2_X4 U32573 ( .A1(n22723), .A2(n22722), .ZN(n22724) );
NAND2_X4 U32574 ( .A1(n20594), .A2(n22724), .ZN(n22737) );
NAND2_X4 U32575 ( .A1(n20630), .A2(n22725), .ZN(n22735) );
NAND2_X4 U32576 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n22863) );
NAND2_X4 U32577 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n22726) );
OR2_X4 U32578 ( .A1(n22726), .A2(n22727), .ZN(n22729) );
NAND2_X4 U32579 ( .A1(n22727), .A2(n22726), .ZN(n22728) );
NAND2_X4 U32580 ( .A1(n22729), .A2(n22728), .ZN(n22731) );
NAND2_X4 U32581 ( .A1(n20627), .A2(n22731), .ZN(n22734) );
NOR2_X4 U32582 ( .A1(n16200), .A2(n20798), .ZN(n22730) );
NOR2_X4 U32583 ( .A1(n20801), .A2(n20675), .ZN(n22872) );
NAND2_X4 U32584 ( .A1(n22730), .A2(n22872), .ZN(n22862) );
NAND2_X4 U32585 ( .A1(n20660), .A2(n22863), .ZN(n22732) );
NAND2_X4 U32586 ( .A1(n20658), .A2(n22732), .ZN(n22733) );
NAND2_X4 U32587 ( .A1(n22734), .A2(n22733), .ZN(n22854) );
NAND2_X4 U32588 ( .A1(n22735), .A2(n22854), .ZN(n22736) );
NAND2_X4 U32589 ( .A1(n22737), .A2(n22736), .ZN(n22846) );
NAND2_X4 U32590 ( .A1(n22738), .A2(n22846), .ZN(n22739) );
NAND2_X4 U32591 ( .A1(n22740), .A2(n22739), .ZN(n22838) );
NAND2_X4 U32592 ( .A1(n22741), .A2(n22838), .ZN(n22742) );
NAND2_X4 U32593 ( .A1(n22743), .A2(n22742), .ZN(n22830) );
NAND2_X4 U32594 ( .A1(n22744), .A2(n22830), .ZN(n22745) );
NAND2_X4 U32595 ( .A1(n22746), .A2(n22745), .ZN(n22822) );
NAND2_X4 U32596 ( .A1(n22747), .A2(n22822), .ZN(n22748) );
NAND2_X4 U32597 ( .A1(n22749), .A2(n22748), .ZN(n22906) );
NAND2_X4 U32598 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n22904) );
OR2_X4 U32599 ( .A1(n22906), .A2(n20403), .ZN(n22751) );
NAND2_X4 U32600 ( .A1(n20403), .A2(n22906), .ZN(n22750) );
NAND2_X4 U32601 ( .A1(n22751), .A2(n22750), .ZN(n22817) );
NAND2_X4 U32602 ( .A1(n20482), .A2(n20519), .ZN(n22757) );
NAND2_X4 U32603 ( .A1(n22753), .A2(n22752), .ZN(n22755) );
NAND2_X4 U32604 ( .A1(n22755), .A2(n22754), .ZN(n22756) );
NAND2_X4 U32605 ( .A1(n22757), .A2(n22756), .ZN(n22914) );
NAND2_X4 U32606 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n22913) );
OR2_X4 U32607 ( .A1(n22914), .A2(n20440), .ZN(n22759) );
NAND2_X4 U32608 ( .A1(n20440), .A2(n22914), .ZN(n22758) );
NAND2_X4 U32609 ( .A1(n22759), .A2(n22758), .ZN(n22814) );
NAND2_X4 U32610 ( .A1(n20520), .A2(n22760), .ZN(n22765) );
NAND2_X4 U32611 ( .A1(n20557), .A2(n22761), .ZN(n22763) );
NAND2_X4 U32612 ( .A1(n22763), .A2(n22762), .ZN(n22764) );
NAND2_X4 U32613 ( .A1(n22765), .A2(n22764), .ZN(n22922) );
NAND2_X4 U32614 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n22920) );
OR2_X4 U32615 ( .A1(n22922), .A2(n20478), .ZN(n22767) );
NAND2_X4 U32616 ( .A1(n20478), .A2(n22922), .ZN(n22766) );
NAND2_X4 U32617 ( .A1(n22767), .A2(n22766), .ZN(n22811) );
NAND2_X4 U32618 ( .A1(n20558), .A2(n20595), .ZN(n22773) );
NAND2_X4 U32619 ( .A1(n22769), .A2(n22768), .ZN(n22771) );
NAND2_X4 U32620 ( .A1(n22771), .A2(n22770), .ZN(n22772) );
NAND2_X4 U32621 ( .A1(n22773), .A2(n22772), .ZN(n22930) );
NAND2_X4 U32622 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n22929) );
OR2_X4 U32623 ( .A1(n22930), .A2(n20516), .ZN(n22775) );
NAND2_X4 U32624 ( .A1(n20516), .A2(n22930), .ZN(n22774) );
NAND2_X4 U32625 ( .A1(n22775), .A2(n22774), .ZN(n22808) );
NAND2_X4 U32626 ( .A1(n20596), .A2(n22776), .ZN(n22781) );
NAND2_X4 U32627 ( .A1(n20628), .A2(n22777), .ZN(n22779) );
NAND2_X4 U32628 ( .A1(n22779), .A2(n22778), .ZN(n22780) );
NAND2_X4 U32629 ( .A1(n22781), .A2(n22780), .ZN(n22938) );
NAND2_X4 U32630 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n22936) );
OR2_X4 U32631 ( .A1(n22938), .A2(n20554), .ZN(n22783) );
NAND2_X4 U32632 ( .A1(n20554), .A2(n22938), .ZN(n22782) );
NAND2_X4 U32633 ( .A1(n22783), .A2(n22782), .ZN(n22805) );
NAND2_X4 U32634 ( .A1(n20629), .A2(n22784), .ZN(n22788) );
NAND2_X4 U32635 ( .A1(n20659), .A2(n22785), .ZN(n22786) );
NAND2_X4 U32636 ( .A1(n20662), .A2(n22786), .ZN(n22787) );
NAND2_X4 U32637 ( .A1(n22788), .A2(n22787), .ZN(n22946) );
NAND2_X4 U32638 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n22945) );
OR2_X4 U32639 ( .A1(n22946), .A2(n20592), .ZN(n22790) );
NAND2_X4 U32640 ( .A1(n20592), .A2(n22946), .ZN(n22789) );
NAND2_X4 U32641 ( .A1(n22790), .A2(n22789), .ZN(n22802) );
NAND2_X4 U32642 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n22953) );
NOR2_X4 U32643 ( .A1(n20683), .A2(n20780), .ZN(n22792) );
NAND2_X4 U32644 ( .A1(n22792), .A2(n22791), .ZN(n22793) );
NAND2_X4 U32645 ( .A1(n20625), .A2(n22793), .ZN(n22795) );
NAND2_X4 U32646 ( .A1(n16329), .A2(n22953), .ZN(n22794) );
NAND2_X4 U32647 ( .A1(n22795), .A2(n22794), .ZN(n22799) );
NAND2_X4 U32648 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n22796) );
NOR2_X4 U32649 ( .A1(n20780), .A2(n20675), .ZN(n22959) );
OR2_X4 U32650 ( .A1(n22796), .A2(n22959), .ZN(n22798) );
NAND2_X4 U32651 ( .A1(n22959), .A2(n22796), .ZN(n22797) );
NAND2_X4 U32652 ( .A1(n22798), .A2(n22797), .ZN(n22952) );
NAND2_X4 U32653 ( .A1(n22799), .A2(n20656), .ZN(n22801) );
OR2_X4 U32654 ( .A1(n20656), .A2(n22799), .ZN(n22800) );
NAND2_X4 U32655 ( .A1(n22801), .A2(n22800), .ZN(n22944) );
NAND2_X4 U32656 ( .A1(n22802), .A2(n20624), .ZN(n22804) );
OR2_X4 U32657 ( .A1(n20624), .A2(n22802), .ZN(n22803) );
NAND2_X4 U32658 ( .A1(n22804), .A2(n22803), .ZN(n22937) );
NAND2_X4 U32659 ( .A1(n22805), .A2(n20591), .ZN(n22807) );
OR2_X4 U32660 ( .A1(n20591), .A2(n22805), .ZN(n22806) );
NAND2_X4 U32661 ( .A1(n22807), .A2(n22806), .ZN(n22928) );
NAND2_X4 U32662 ( .A1(n22808), .A2(n20553), .ZN(n22810) );
OR2_X4 U32663 ( .A1(n20553), .A2(n22808), .ZN(n22809) );
NAND2_X4 U32664 ( .A1(n22810), .A2(n22809), .ZN(n22921) );
NAND2_X4 U32665 ( .A1(n22811), .A2(n20515), .ZN(n22813) );
OR2_X4 U32666 ( .A1(n20515), .A2(n22811), .ZN(n22812) );
NAND2_X4 U32667 ( .A1(n22813), .A2(n22812), .ZN(n22912) );
NAND2_X4 U32668 ( .A1(n22814), .A2(n20477), .ZN(n22816) );
OR2_X4 U32669 ( .A1(n20477), .A2(n22814), .ZN(n22815) );
NAND2_X4 U32670 ( .A1(n22816), .A2(n22815), .ZN(n22905) );
NAND2_X4 U32671 ( .A1(n22817), .A2(n20439), .ZN(n22819) );
OR2_X4 U32672 ( .A1(n20439), .A2(n22817), .ZN(n22818) );
NAND2_X4 U32673 ( .A1(n22819), .A2(n22818), .ZN(n22820) );
NAND2_X4 U32674 ( .A1(n20364), .A2(n22820), .ZN(n22901) );
NAND2_X4 U32675 ( .A1(n20402), .A2(n22821), .ZN(n22899) );
NAND2_X4 U32676 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n22828) );
OR2_X4 U32677 ( .A1(n22822), .A2(n20442), .ZN(n22824) );
NAND2_X4 U32678 ( .A1(n20442), .A2(n22822), .ZN(n22823) );
NAND2_X4 U32679 ( .A1(n22824), .A2(n22823), .ZN(n22825) );
NAND2_X4 U32680 ( .A1(n22825), .A2(n20481), .ZN(n22827) );
OR2_X4 U32681 ( .A1(n20481), .A2(n22825), .ZN(n22826) );
NAND2_X4 U32682 ( .A1(n22827), .A2(n22826), .ZN(n22829) );
NAND2_X4 U32683 ( .A1(n20401), .A2(n20441), .ZN(n22898) );
NAND2_X4 U32684 ( .A1(n22829), .A2(n22828), .ZN(n22896) );
NAND2_X4 U32685 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n22837) );
OR2_X4 U32686 ( .A1(n22830), .A2(n20480), .ZN(n22832) );
NAND2_X4 U32687 ( .A1(n20480), .A2(n22830), .ZN(n22831) );
NAND2_X4 U32688 ( .A1(n22832), .A2(n22831), .ZN(n22833) );
NAND2_X4 U32689 ( .A1(n22833), .A2(n20521), .ZN(n22835) );
OR2_X4 U32690 ( .A1(n20521), .A2(n22833), .ZN(n22834) );
NAND2_X4 U32691 ( .A1(n22835), .A2(n22834), .ZN(n22836) );
NAND2_X4 U32692 ( .A1(n20438), .A2(n22836), .ZN(n22895) );
NAND2_X4 U32693 ( .A1(n20479), .A2(n22837), .ZN(n22893) );
NAND2_X4 U32694 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n22844) );
OR2_X4 U32695 ( .A1(n22838), .A2(n20518), .ZN(n22840) );
NAND2_X4 U32696 ( .A1(n20518), .A2(n22838), .ZN(n22839) );
NAND2_X4 U32697 ( .A1(n22840), .A2(n22839), .ZN(n22841) );
NAND2_X4 U32698 ( .A1(n22841), .A2(n20559), .ZN(n22843) );
OR2_X4 U32699 ( .A1(n20559), .A2(n22841), .ZN(n22842) );
NAND2_X4 U32700 ( .A1(n22843), .A2(n22842), .ZN(n22845) );
NAND2_X4 U32701 ( .A1(n20476), .A2(n20517), .ZN(n22892) );
NAND2_X4 U32702 ( .A1(n22845), .A2(n22844), .ZN(n22890) );
NAND2_X4 U32703 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n22853) );
OR2_X4 U32704 ( .A1(n22846), .A2(n20556), .ZN(n22848) );
NAND2_X4 U32705 ( .A1(n20556), .A2(n22846), .ZN(n22847) );
NAND2_X4 U32706 ( .A1(n22848), .A2(n22847), .ZN(n22849) );
NAND2_X4 U32707 ( .A1(n22849), .A2(n20597), .ZN(n22851) );
OR2_X4 U32708 ( .A1(n20597), .A2(n22849), .ZN(n22850) );
NAND2_X4 U32709 ( .A1(n22851), .A2(n22850), .ZN(n22852) );
NAND2_X4 U32710 ( .A1(n20514), .A2(n22852), .ZN(n22889) );
NAND2_X4 U32711 ( .A1(n20555), .A2(n22853), .ZN(n22887) );
NAND2_X4 U32712 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n22860) );
OR2_X4 U32713 ( .A1(n22854), .A2(n20594), .ZN(n22856) );
NAND2_X4 U32714 ( .A1(n20594), .A2(n22854), .ZN(n22855) );
NAND2_X4 U32715 ( .A1(n22856), .A2(n22855), .ZN(n22857) );
NAND2_X4 U32716 ( .A1(n22857), .A2(n20630), .ZN(n22859) );
OR2_X4 U32717 ( .A1(n20630), .A2(n22857), .ZN(n22858) );
NAND2_X4 U32718 ( .A1(n22859), .A2(n22858), .ZN(n22861) );
NAND2_X4 U32719 ( .A1(n20552), .A2(n20593), .ZN(n22886) );
NAND2_X4 U32720 ( .A1(n22861), .A2(n22860), .ZN(n22884) );
NAND2_X4 U32721 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n22870) );
NAND2_X4 U32722 ( .A1(n20627), .A2(n22862), .ZN(n22865) );
NAND2_X4 U32723 ( .A1(n20658), .A2(n22863), .ZN(n22864) );
NAND2_X4 U32724 ( .A1(n22865), .A2(n22864), .ZN(n22866) );
NAND2_X4 U32725 ( .A1(n22866), .A2(n20660), .ZN(n22868) );
OR2_X4 U32726 ( .A1(n20660), .A2(n22866), .ZN(n22867) );
NAND2_X4 U32727 ( .A1(n22868), .A2(n22867), .ZN(n22869) );
NAND2_X4 U32728 ( .A1(n20590), .A2(n22869), .ZN(n22883) );
NAND2_X4 U32729 ( .A1(n20626), .A2(n22870), .ZN(n22881) );
NAND2_X4 U32730 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n23037) );
NAND2_X4 U32731 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n22871) );
OR2_X4 U32732 ( .A1(n22871), .A2(n22872), .ZN(n22874) );
NAND2_X4 U32733 ( .A1(n22872), .A2(n22871), .ZN(n22873) );
NAND2_X4 U32734 ( .A1(n22874), .A2(n22873), .ZN(n22877) );
NAND2_X4 U32735 ( .A1(n20623), .A2(n22877), .ZN(n22880) );
NOR2_X4 U32736 ( .A1(n16200), .A2(n20801), .ZN(n22876) );
NAND2_X4 U32737 ( .A1(n22876), .A2(n22875), .ZN(n23036) );
NAND2_X4 U32738 ( .A1(n20657), .A2(n23037), .ZN(n22878) );
NAND2_X4 U32739 ( .A1(n20670), .A2(n22878), .ZN(n22879) );
NAND2_X4 U32740 ( .A1(n22880), .A2(n22879), .ZN(n23030) );
NAND2_X4 U32741 ( .A1(n22881), .A2(n23030), .ZN(n22882) );
NAND2_X4 U32742 ( .A1(n22883), .A2(n22882), .ZN(n23024) );
NAND2_X4 U32743 ( .A1(n22884), .A2(n23024), .ZN(n22885) );
NAND2_X4 U32744 ( .A1(n22886), .A2(n22885), .ZN(n23018) );
NAND2_X4 U32745 ( .A1(n22887), .A2(n23018), .ZN(n22888) );
NAND2_X4 U32746 ( .A1(n22889), .A2(n22888), .ZN(n23012) );
NAND2_X4 U32747 ( .A1(n22890), .A2(n23012), .ZN(n22891) );
NAND2_X4 U32748 ( .A1(n22892), .A2(n22891), .ZN(n23006) );
NAND2_X4 U32749 ( .A1(n22893), .A2(n23006), .ZN(n22894) );
NAND2_X4 U32750 ( .A1(n22895), .A2(n22894), .ZN(n23000) );
NAND2_X4 U32751 ( .A1(n22896), .A2(n23000), .ZN(n22897) );
NAND2_X4 U32752 ( .A1(n22898), .A2(n22897), .ZN(n22994) );
NAND2_X4 U32753 ( .A1(n22899), .A2(n22994), .ZN(n22900) );
NAND2_X4 U32754 ( .A1(n22901), .A2(n22900), .ZN(n23090) );
NAND2_X4 U32755 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n23088) );
OR2_X4 U32756 ( .A1(n23090), .A2(n20325), .ZN(n22903) );
NAND2_X4 U32757 ( .A1(n20325), .A2(n23090), .ZN(n22902) );
NAND2_X4 U32758 ( .A1(n22903), .A2(n22902), .ZN(n22991) );
NAND2_X4 U32759 ( .A1(n20403), .A2(n20439), .ZN(n22909) );
NAND2_X4 U32760 ( .A1(n22905), .A2(n22904), .ZN(n22907) );
NAND2_X4 U32761 ( .A1(n22907), .A2(n22906), .ZN(n22908) );
NAND2_X4 U32762 ( .A1(n22909), .A2(n22908), .ZN(n23098) );
NAND2_X4 U32763 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n23097) );
OR2_X4 U32764 ( .A1(n23098), .A2(n20362), .ZN(n22911) );
NAND2_X4 U32765 ( .A1(n20362), .A2(n23098), .ZN(n22910) );
NAND2_X4 U32766 ( .A1(n22911), .A2(n22910), .ZN(n22988) );
NAND2_X4 U32767 ( .A1(n20440), .A2(n22912), .ZN(n22917) );
NAND2_X4 U32768 ( .A1(n20477), .A2(n22913), .ZN(n22915) );
NAND2_X4 U32769 ( .A1(n22915), .A2(n22914), .ZN(n22916) );
NAND2_X4 U32770 ( .A1(n22917), .A2(n22916), .ZN(n23106) );
NAND2_X4 U32771 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n23104) );
OR2_X4 U32772 ( .A1(n23106), .A2(n20399), .ZN(n22919) );
NAND2_X4 U32773 ( .A1(n20399), .A2(n23106), .ZN(n22918) );
NAND2_X4 U32774 ( .A1(n22919), .A2(n22918), .ZN(n22985) );
NAND2_X4 U32775 ( .A1(n20478), .A2(n20515), .ZN(n22925) );
NAND2_X4 U32776 ( .A1(n22921), .A2(n22920), .ZN(n22923) );
NAND2_X4 U32777 ( .A1(n22923), .A2(n22922), .ZN(n22924) );
NAND2_X4 U32778 ( .A1(n22925), .A2(n22924), .ZN(n23114) );
NAND2_X4 U32779 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n23113) );
OR2_X4 U32780 ( .A1(n23114), .A2(n20436), .ZN(n22927) );
NAND2_X4 U32781 ( .A1(n20436), .A2(n23114), .ZN(n22926) );
NAND2_X4 U32782 ( .A1(n22927), .A2(n22926), .ZN(n22982) );
NAND2_X4 U32783 ( .A1(n20516), .A2(n22928), .ZN(n22933) );
NAND2_X4 U32784 ( .A1(n20553), .A2(n22929), .ZN(n22931) );
NAND2_X4 U32785 ( .A1(n22931), .A2(n22930), .ZN(n22932) );
NAND2_X4 U32786 ( .A1(n22933), .A2(n22932), .ZN(n23122) );
NAND2_X4 U32787 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n23120) );
OR2_X4 U32788 ( .A1(n23122), .A2(n20474), .ZN(n22935) );
NAND2_X4 U32789 ( .A1(n20474), .A2(n23122), .ZN(n22934) );
NAND2_X4 U32790 ( .A1(n22935), .A2(n22934), .ZN(n22979) );
NAND2_X4 U32791 ( .A1(n20554), .A2(n20591), .ZN(n22941) );
NAND2_X4 U32792 ( .A1(n22937), .A2(n22936), .ZN(n22939) );
NAND2_X4 U32793 ( .A1(n22939), .A2(n22938), .ZN(n22940) );
NAND2_X4 U32794 ( .A1(n22941), .A2(n22940), .ZN(n23130) );
NAND2_X4 U32795 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n23129) );
OR2_X4 U32796 ( .A1(n23130), .A2(n20512), .ZN(n22943) );
NAND2_X4 U32797 ( .A1(n20512), .A2(n23130), .ZN(n22942) );
NAND2_X4 U32798 ( .A1(n22943), .A2(n22942), .ZN(n22976) );
NAND2_X4 U32799 ( .A1(n20592), .A2(n22944), .ZN(n22949) );
NAND2_X4 U32800 ( .A1(n20624), .A2(n22945), .ZN(n22947) );
NAND2_X4 U32801 ( .A1(n22947), .A2(n22946), .ZN(n22948) );
NAND2_X4 U32802 ( .A1(n22949), .A2(n22948), .ZN(n23138) );
NAND2_X4 U32803 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n23136) );
OR2_X4 U32804 ( .A1(n23138), .A2(n20550), .ZN(n22951) );
NAND2_X4 U32805 ( .A1(n20550), .A2(n23138), .ZN(n22950) );
NAND2_X4 U32806 ( .A1(n22951), .A2(n22950), .ZN(n22973) );
NAND2_X4 U32807 ( .A1(n20625), .A2(n22952), .ZN(n22956) );
NAND2_X4 U32808 ( .A1(n20656), .A2(n22953), .ZN(n22954) );
NAND2_X4 U32809 ( .A1(n16329), .A2(n22954), .ZN(n22955) );
NAND2_X4 U32810 ( .A1(n22956), .A2(n22955), .ZN(n23146) );
NAND2_X4 U32811 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n23145) );
OR2_X4 U32812 ( .A1(n23146), .A2(n20588), .ZN(n22958) );
NAND2_X4 U32813 ( .A1(n20588), .A2(n23146), .ZN(n22957) );
NAND2_X4 U32814 ( .A1(n22958), .A2(n22957), .ZN(n22970) );
NAND2_X4 U32815 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n23153) );
NOR2_X4 U32816 ( .A1(n20683), .A2(n20777), .ZN(n22960) );
NAND2_X4 U32817 ( .A1(n22960), .A2(n22959), .ZN(n22961) );
NAND2_X4 U32818 ( .A1(n20621), .A2(n22961), .ZN(n22963) );
NAND2_X4 U32819 ( .A1(n16328), .A2(n23153), .ZN(n22962) );
NAND2_X4 U32820 ( .A1(n22963), .A2(n22962), .ZN(n22967) );
NAND2_X4 U32821 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n22964) );
NOR2_X4 U32822 ( .A1(n20777), .A2(n20675), .ZN(n23159) );
OR2_X4 U32823 ( .A1(n22964), .A2(n23159), .ZN(n22966) );
NAND2_X4 U32824 ( .A1(n23159), .A2(n22964), .ZN(n22965) );
NAND2_X4 U32825 ( .A1(n22966), .A2(n22965), .ZN(n23152) );
NAND2_X4 U32826 ( .A1(n22967), .A2(n20655), .ZN(n22969) );
OR2_X4 U32827 ( .A1(n20655), .A2(n22967), .ZN(n22968) );
NAND2_X4 U32828 ( .A1(n22969), .A2(n22968), .ZN(n23144) );
NAND2_X4 U32829 ( .A1(n22970), .A2(n20620), .ZN(n22972) );
OR2_X4 U32830 ( .A1(n20620), .A2(n22970), .ZN(n22971) );
NAND2_X4 U32831 ( .A1(n22972), .A2(n22971), .ZN(n23137) );
NAND2_X4 U32832 ( .A1(n22973), .A2(n20587), .ZN(n22975) );
OR2_X4 U32833 ( .A1(n20587), .A2(n22973), .ZN(n22974) );
NAND2_X4 U32834 ( .A1(n22975), .A2(n22974), .ZN(n23128) );
NAND2_X4 U32835 ( .A1(n22976), .A2(n20549), .ZN(n22978) );
OR2_X4 U32836 ( .A1(n20549), .A2(n22976), .ZN(n22977) );
NAND2_X4 U32837 ( .A1(n22978), .A2(n22977), .ZN(n23121) );
NAND2_X4 U32838 ( .A1(n22979), .A2(n20511), .ZN(n22981) );
OR2_X4 U32839 ( .A1(n20511), .A2(n22979), .ZN(n22980) );
NAND2_X4 U32840 ( .A1(n22981), .A2(n22980), .ZN(n23112) );
NAND2_X4 U32841 ( .A1(n22982), .A2(n16333), .ZN(n22984) );
OR2_X4 U32842 ( .A1(n16333), .A2(n22982), .ZN(n22983) );
NAND2_X4 U32843 ( .A1(n22984), .A2(n22983), .ZN(n23105) );
NAND2_X4 U32844 ( .A1(n22985), .A2(n20435), .ZN(n22987) );
OR2_X4 U32845 ( .A1(n20435), .A2(n22985), .ZN(n22986) );
NAND2_X4 U32846 ( .A1(n22987), .A2(n22986), .ZN(n23096) );
NAND2_X4 U32847 ( .A1(n22988), .A2(n20398), .ZN(n22990) );
OR2_X4 U32848 ( .A1(n20398), .A2(n22988), .ZN(n22989) );
NAND2_X4 U32849 ( .A1(n22990), .A2(n22989), .ZN(n23089) );
NAND2_X4 U32850 ( .A1(n22991), .A2(n20361), .ZN(n22993) );
OR2_X4 U32851 ( .A1(n20361), .A2(n22991), .ZN(n22992) );
NAND2_X4 U32852 ( .A1(n22993), .A2(n22992), .ZN(n23081) );
OR2_X4 U32853 ( .A1(n22994), .A2(n20364), .ZN(n22996) );
NAND2_X4 U32854 ( .A1(n20364), .A2(n22994), .ZN(n22995) );
NAND2_X4 U32855 ( .A1(n22996), .A2(n22995), .ZN(n22997) );
NAND2_X4 U32856 ( .A1(n22997), .A2(n20402), .ZN(n22999) );
OR2_X4 U32857 ( .A1(n20402), .A2(n22997), .ZN(n22998) );
NAND2_X4 U32858 ( .A1(n22999), .A2(n22998), .ZN(n23077) );
OR2_X4 U32859 ( .A1(n23000), .A2(n20401), .ZN(n23002) );
NAND2_X4 U32860 ( .A1(n20401), .A2(n23000), .ZN(n23001) );
NAND2_X4 U32861 ( .A1(n23002), .A2(n23001), .ZN(n23003) );
NAND2_X4 U32862 ( .A1(n23003), .A2(n20441), .ZN(n23005) );
OR2_X4 U32863 ( .A1(n20441), .A2(n23003), .ZN(n23004) );
NAND2_X4 U32864 ( .A1(n23005), .A2(n23004), .ZN(n23073) );
OR2_X4 U32865 ( .A1(n23006), .A2(n20438), .ZN(n23008) );
NAND2_X4 U32866 ( .A1(n20438), .A2(n23006), .ZN(n23007) );
NAND2_X4 U32867 ( .A1(n23008), .A2(n23007), .ZN(n23009) );
NAND2_X4 U32868 ( .A1(n23009), .A2(n20479), .ZN(n23011) );
OR2_X4 U32869 ( .A1(n20479), .A2(n23009), .ZN(n23010) );
NAND2_X4 U32870 ( .A1(n23011), .A2(n23010), .ZN(n23069) );
OR2_X4 U32871 ( .A1(n23012), .A2(n20476), .ZN(n23014) );
NAND2_X4 U32872 ( .A1(n20476), .A2(n23012), .ZN(n23013) );
NAND2_X4 U32873 ( .A1(n23014), .A2(n23013), .ZN(n23015) );
NAND2_X4 U32874 ( .A1(n23015), .A2(n20517), .ZN(n23017) );
OR2_X4 U32875 ( .A1(n20517), .A2(n23015), .ZN(n23016) );
NAND2_X4 U32876 ( .A1(n23017), .A2(n23016), .ZN(n23065) );
OR2_X4 U32877 ( .A1(n23018), .A2(n20514), .ZN(n23020) );
NAND2_X4 U32878 ( .A1(n20514), .A2(n23018), .ZN(n23019) );
NAND2_X4 U32879 ( .A1(n23020), .A2(n23019), .ZN(n23021) );
NAND2_X4 U32880 ( .A1(n23021), .A2(n20555), .ZN(n23023) );
OR2_X4 U32881 ( .A1(n20555), .A2(n23021), .ZN(n23022) );
NAND2_X4 U32882 ( .A1(n23023), .A2(n23022), .ZN(n23061) );
OR2_X4 U32883 ( .A1(n23024), .A2(n20552), .ZN(n23026) );
NAND2_X4 U32884 ( .A1(n20552), .A2(n23024), .ZN(n23025) );
NAND2_X4 U32885 ( .A1(n23026), .A2(n23025), .ZN(n23027) );
NAND2_X4 U32886 ( .A1(n23027), .A2(n20593), .ZN(n23029) );
OR2_X4 U32887 ( .A1(n20593), .A2(n23027), .ZN(n23028) );
NAND2_X4 U32888 ( .A1(n23029), .A2(n23028), .ZN(n23057) );
OR2_X4 U32889 ( .A1(n23030), .A2(n20590), .ZN(n23032) );
NAND2_X4 U32890 ( .A1(n20590), .A2(n23030), .ZN(n23031) );
NAND2_X4 U32891 ( .A1(n23032), .A2(n23031), .ZN(n23033) );
NAND2_X4 U32892 ( .A1(n23033), .A2(n20626), .ZN(n23035) );
OR2_X4 U32893 ( .A1(n20626), .A2(n23033), .ZN(n23034) );
NAND2_X4 U32894 ( .A1(n23035), .A2(n23034), .ZN(n23053) );
NAND2_X4 U32895 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n23044) );
NAND2_X4 U32896 ( .A1(n20623), .A2(n23036), .ZN(n23039) );
NAND2_X4 U32897 ( .A1(n20670), .A2(n23037), .ZN(n23038) );
NAND2_X4 U32898 ( .A1(n23039), .A2(n23038), .ZN(n23040) );
NAND2_X4 U32899 ( .A1(n23040), .A2(n20657), .ZN(n23042) );
OR2_X4 U32900 ( .A1(n20657), .A2(n23040), .ZN(n23041) );
NAND2_X4 U32901 ( .A1(n23042), .A2(n23041), .ZN(n23043) );
NAND2_X4 U32902 ( .A1(n20586), .A2(n23043), .ZN(n23052) );
NAND2_X4 U32903 ( .A1(n20622), .A2(n23044), .ZN(n23050) );
NAND2_X4 U32904 ( .A1(n20674), .A2(n23045), .ZN(n23049) );
NAND2_X4 U32905 ( .A1(n20671), .A2(n23046), .ZN(n23047) );
NAND2_X4 U32906 ( .A1(n20640), .A2(n23047), .ZN(n23048) );
NAND2_X4 U32907 ( .A1(n23049), .A2(n23048), .ZN(n24524) );
NAND2_X4 U32908 ( .A1(n23050), .A2(n24524), .ZN(n23051) );
NAND2_X4 U32909 ( .A1(n23052), .A2(n23051), .ZN(n25185) );
NAND2_X4 U32910 ( .A1(n20589), .A2(n25185), .ZN(n23056) );
NAND2_X4 U32911 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n25184) );
NAND2_X4 U32912 ( .A1(n20583), .A2(n23053), .ZN(n23054) );
NAND2_X4 U32913 ( .A1(n20548), .A2(n23054), .ZN(n23055) );
NAND2_X4 U32914 ( .A1(n23056), .A2(n23055), .ZN(n25195) );
NAND2_X4 U32915 ( .A1(n23057), .A2(n25195), .ZN(n23060) );
NAND2_X4 U32916 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n25194) );
NAND2_X4 U32917 ( .A1(n20547), .A2(n20551), .ZN(n23058) );
NAND2_X4 U32918 ( .A1(n20510), .A2(n23058), .ZN(n23059) );
NAND2_X4 U32919 ( .A1(n23060), .A2(n23059), .ZN(n25202) );
NAND2_X4 U32920 ( .A1(n20513), .A2(n25202), .ZN(n23064) );
NAND2_X4 U32921 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n25201) );
NAND2_X4 U32922 ( .A1(n20509), .A2(n23061), .ZN(n23062) );
NAND2_X4 U32923 ( .A1(n20472), .A2(n23062), .ZN(n23063) );
NAND2_X4 U32924 ( .A1(n23064), .A2(n23063), .ZN(n25209) );
NAND2_X4 U32925 ( .A1(n23065), .A2(n25209), .ZN(n23068) );
NAND2_X4 U32926 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n25208) );
NAND2_X4 U32927 ( .A1(n20471), .A2(n20475), .ZN(n23066) );
NAND2_X4 U32928 ( .A1(n20434), .A2(n23066), .ZN(n23067) );
NAND2_X4 U32929 ( .A1(n23068), .A2(n23067), .ZN(n25216) );
NAND2_X4 U32930 ( .A1(n20437), .A2(n25216), .ZN(n23072) );
NAND2_X4 U32931 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n25215) );
NAND2_X4 U32932 ( .A1(n20433), .A2(n23069), .ZN(n23070) );
NAND2_X4 U32933 ( .A1(n20397), .A2(n23070), .ZN(n23071) );
NAND2_X4 U32934 ( .A1(n23072), .A2(n23071), .ZN(n25223) );
NAND2_X4 U32935 ( .A1(n23073), .A2(n25223), .ZN(n23076) );
NAND2_X4 U32936 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n25222) );
NAND2_X4 U32937 ( .A1(n20396), .A2(n20400), .ZN(n23074) );
NAND2_X4 U32938 ( .A1(n20360), .A2(n23074), .ZN(n23075) );
NAND2_X4 U32939 ( .A1(n23076), .A2(n23075), .ZN(n25230) );
NAND2_X4 U32940 ( .A1(n20363), .A2(n25230), .ZN(n23080) );
NAND2_X4 U32941 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n25229) );
NAND2_X4 U32942 ( .A1(n20359), .A2(n23077), .ZN(n23078) );
NAND2_X4 U32943 ( .A1(n20323), .A2(n23078), .ZN(n23079) );
NAND2_X4 U32944 ( .A1(n23080), .A2(n23079), .ZN(n25237) );
NAND2_X4 U32945 ( .A1(n23081), .A2(n25237), .ZN(n23084) );
NAND2_X4 U32946 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n25236) );
NAND2_X4 U32947 ( .A1(n20322), .A2(n20324), .ZN(n23082) );
NAND2_X4 U32948 ( .A1(n20286), .A2(n23082), .ZN(n23083) );
NAND2_X4 U32949 ( .A1(n23084), .A2(n23083), .ZN(n23200) );
NAND2_X4 U32950 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n23085) );
NAND2_X4 U32951 ( .A1(n20285), .A2(n23085), .ZN(n23087) );
NAND2_X4 U32952 ( .A1(n20247), .A2(n23200), .ZN(n23086) );
NAND2_X4 U32953 ( .A1(n23087), .A2(n23086), .ZN(n23197) );
NAND2_X4 U32954 ( .A1(n20325), .A2(n20361), .ZN(n23093) );
NAND2_X4 U32955 ( .A1(n23089), .A2(n23088), .ZN(n23091) );
NAND2_X4 U32956 ( .A1(n23091), .A2(n23090), .ZN(n23092) );
NAND2_X4 U32957 ( .A1(n23093), .A2(n23092), .ZN(n23209) );
NAND2_X4 U32958 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n23208) );
OR2_X4 U32959 ( .A1(n23209), .A2(n20282), .ZN(n23095) );
NAND2_X4 U32960 ( .A1(n20282), .A2(n23209), .ZN(n23094) );
NAND2_X4 U32961 ( .A1(n23095), .A2(n23094), .ZN(n23194) );
NAND2_X4 U32962 ( .A1(n20362), .A2(n23096), .ZN(n23101) );
NAND2_X4 U32963 ( .A1(n20398), .A2(n23097), .ZN(n23099) );
NAND2_X4 U32964 ( .A1(n23099), .A2(n23098), .ZN(n23100) );
NAND2_X4 U32965 ( .A1(n23101), .A2(n23100), .ZN(n23217) );
NAND2_X4 U32966 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n23215) );
OR2_X4 U32967 ( .A1(n23217), .A2(n20319), .ZN(n23103) );
NAND2_X4 U32968 ( .A1(n20319), .A2(n23217), .ZN(n23102) );
NAND2_X4 U32969 ( .A1(n23103), .A2(n23102), .ZN(n23191) );
NAND2_X4 U32970 ( .A1(n20399), .A2(n20435), .ZN(n23109) );
NAND2_X4 U32971 ( .A1(n23105), .A2(n23104), .ZN(n23107) );
NAND2_X4 U32972 ( .A1(n23107), .A2(n23106), .ZN(n23108) );
NAND2_X4 U32973 ( .A1(n23109), .A2(n23108), .ZN(n23225) );
NAND2_X4 U32974 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n23224) );
OR2_X4 U32975 ( .A1(n23225), .A2(n20356), .ZN(n23111) );
NAND2_X4 U32976 ( .A1(n20356), .A2(n23225), .ZN(n23110) );
NAND2_X4 U32977 ( .A1(n23111), .A2(n23110), .ZN(n23188) );
NAND2_X4 U32978 ( .A1(n20436), .A2(n23112), .ZN(n23117) );
NAND2_X4 U32979 ( .A1(n20473), .A2(n23113), .ZN(n23115) );
NAND2_X4 U32980 ( .A1(n23115), .A2(n23114), .ZN(n23116) );
NAND2_X4 U32981 ( .A1(n23117), .A2(n23116), .ZN(n23233) );
NAND2_X4 U32982 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n23231) );
OR2_X4 U32983 ( .A1(n23233), .A2(n20393), .ZN(n23119) );
NAND2_X4 U32984 ( .A1(n20393), .A2(n23233), .ZN(n23118) );
NAND2_X4 U32985 ( .A1(n23119), .A2(n23118), .ZN(n23185) );
NAND2_X4 U32986 ( .A1(n20474), .A2(n20511), .ZN(n23125) );
NAND2_X4 U32987 ( .A1(n23121), .A2(n23120), .ZN(n23123) );
NAND2_X4 U32988 ( .A1(n23123), .A2(n23122), .ZN(n23124) );
NAND2_X4 U32989 ( .A1(n23125), .A2(n23124), .ZN(n23241) );
NAND2_X4 U32990 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n23240) );
OR2_X4 U32991 ( .A1(n23241), .A2(n20430), .ZN(n23127) );
NAND2_X4 U32992 ( .A1(n20430), .A2(n23241), .ZN(n23126) );
NAND2_X4 U32993 ( .A1(n23127), .A2(n23126), .ZN(n23182) );
NAND2_X4 U32994 ( .A1(n20512), .A2(n23128), .ZN(n23133) );
NAND2_X4 U32995 ( .A1(n20549), .A2(n23129), .ZN(n23131) );
NAND2_X4 U32996 ( .A1(n23131), .A2(n23130), .ZN(n23132) );
NAND2_X4 U32997 ( .A1(n23133), .A2(n23132), .ZN(n23249) );
NAND2_X4 U32998 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n23247) );
OR2_X4 U32999 ( .A1(n23249), .A2(n20468), .ZN(n23135) );
NAND2_X4 U33000 ( .A1(n20468), .A2(n23249), .ZN(n23134) );
NAND2_X4 U33001 ( .A1(n23135), .A2(n23134), .ZN(n23179) );
NAND2_X4 U33002 ( .A1(n20550), .A2(n20587), .ZN(n23141) );
NAND2_X4 U33003 ( .A1(n23137), .A2(n23136), .ZN(n23139) );
NAND2_X4 U33004 ( .A1(n23139), .A2(n23138), .ZN(n23140) );
NAND2_X4 U33005 ( .A1(n23141), .A2(n23140), .ZN(n23257) );
NAND2_X4 U33006 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n23256) );
OR2_X4 U33007 ( .A1(n23257), .A2(n20506), .ZN(n23143) );
NAND2_X4 U33008 ( .A1(n20506), .A2(n23257), .ZN(n23142) );
NAND2_X4 U33009 ( .A1(n23143), .A2(n23142), .ZN(n23176) );
NAND2_X4 U33010 ( .A1(n20588), .A2(n23144), .ZN(n23149) );
NAND2_X4 U33011 ( .A1(n20620), .A2(n23145), .ZN(n23147) );
NAND2_X4 U33012 ( .A1(n23147), .A2(n23146), .ZN(n23148) );
NAND2_X4 U33013 ( .A1(n23149), .A2(n23148), .ZN(n23265) );
NAND2_X4 U33014 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n23263) );
OR2_X4 U33015 ( .A1(n23265), .A2(n20544), .ZN(n23151) );
NAND2_X4 U33016 ( .A1(n20544), .A2(n23265), .ZN(n23150) );
NAND2_X4 U33017 ( .A1(n23151), .A2(n23150), .ZN(n23173) );
NAND2_X4 U33018 ( .A1(n20621), .A2(n23152), .ZN(n23156) );
NAND2_X4 U33019 ( .A1(n20655), .A2(n23153), .ZN(n23154) );
NAND2_X4 U33020 ( .A1(n16328), .A2(n23154), .ZN(n23155) );
NAND2_X4 U33021 ( .A1(n23156), .A2(n23155), .ZN(n23273) );
NAND2_X4 U33022 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n23272) );
OR2_X4 U33023 ( .A1(n23273), .A2(n20582), .ZN(n23158) );
NAND2_X4 U33024 ( .A1(n20582), .A2(n23273), .ZN(n23157) );
NAND2_X4 U33025 ( .A1(n23158), .A2(n23157), .ZN(n23170) );
NAND2_X4 U33026 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n23280) );
NOR2_X4 U33027 ( .A1(n16200), .A2(n20774), .ZN(n23160) );
NAND2_X4 U33028 ( .A1(n23160), .A2(n23159), .ZN(n23161) );
NAND2_X4 U33029 ( .A1(n20619), .A2(n23161), .ZN(n23163) );
NAND2_X4 U33030 ( .A1(n20654), .A2(n23280), .ZN(n23162) );
NAND2_X4 U33031 ( .A1(n23163), .A2(n23162), .ZN(n23167) );
NAND2_X4 U33032 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n23164) );
NOR2_X4 U33033 ( .A1(n20774), .A2(n20675), .ZN(n23286) );
OR2_X4 U33034 ( .A1(n23164), .A2(n23286), .ZN(n23166) );
NAND2_X4 U33035 ( .A1(n23286), .A2(n23164), .ZN(n23165) );
NAND2_X4 U33036 ( .A1(n23166), .A2(n23165), .ZN(n23279) );
NAND2_X4 U33037 ( .A1(n23167), .A2(n20653), .ZN(n23169) );
OR2_X4 U33038 ( .A1(n20653), .A2(n23167), .ZN(n23168) );
NAND2_X4 U33039 ( .A1(n23169), .A2(n23168), .ZN(n23271) );
NAND2_X4 U33040 ( .A1(n23170), .A2(n20618), .ZN(n23172) );
OR2_X4 U33041 ( .A1(n20618), .A2(n23170), .ZN(n23171) );
NAND2_X4 U33042 ( .A1(n23172), .A2(n23171), .ZN(n23264) );
NAND2_X4 U33043 ( .A1(n23173), .A2(n20581), .ZN(n23175) );
OR2_X4 U33044 ( .A1(n20581), .A2(n23173), .ZN(n23174) );
NAND2_X4 U33045 ( .A1(n23175), .A2(n23174), .ZN(n23255) );
NAND2_X4 U33046 ( .A1(n23176), .A2(n20543), .ZN(n23178) );
OR2_X4 U33047 ( .A1(n20543), .A2(n23176), .ZN(n23177) );
NAND2_X4 U33048 ( .A1(n23178), .A2(n23177), .ZN(n23248) );
NAND2_X4 U33049 ( .A1(n23179), .A2(n20505), .ZN(n23181) );
OR2_X4 U33050 ( .A1(n20505), .A2(n23179), .ZN(n23180) );
NAND2_X4 U33051 ( .A1(n23181), .A2(n23180), .ZN(n23239) );
NAND2_X4 U33052 ( .A1(n23182), .A2(n20467), .ZN(n23184) );
OR2_X4 U33053 ( .A1(n20467), .A2(n23182), .ZN(n23183) );
NAND2_X4 U33054 ( .A1(n23184), .A2(n23183), .ZN(n23232) );
NAND2_X4 U33055 ( .A1(n23185), .A2(n20429), .ZN(n23187) );
OR2_X4 U33056 ( .A1(n20429), .A2(n23185), .ZN(n23186) );
NAND2_X4 U33057 ( .A1(n23187), .A2(n23186), .ZN(n23223) );
NAND2_X4 U33058 ( .A1(n23188), .A2(n16332), .ZN(n23190) );
OR2_X4 U33059 ( .A1(n16332), .A2(n23188), .ZN(n23189) );
NAND2_X4 U33060 ( .A1(n23190), .A2(n23189), .ZN(n23216) );
NAND2_X4 U33061 ( .A1(n23191), .A2(n20355), .ZN(n23193) );
OR2_X4 U33062 ( .A1(n20355), .A2(n23191), .ZN(n23192) );
NAND2_X4 U33063 ( .A1(n23193), .A2(n23192), .ZN(n23207) );
NAND2_X4 U33064 ( .A1(n23194), .A2(n20318), .ZN(n23196) );
OR2_X4 U33065 ( .A1(n20318), .A2(n23194), .ZN(n23195) );
NAND2_X4 U33066 ( .A1(n23196), .A2(n23195), .ZN(n23201) );
NAND2_X4 U33067 ( .A1(n23197), .A2(n20281), .ZN(n23199) );
OR2_X4 U33068 ( .A1(n20281), .A2(n23197), .ZN(n23198) );
NAND2_X4 U33069 ( .A1(n23199), .A2(n23198), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N47) );
NAND2_X4 U33070 ( .A1(n20281), .A2(n23200), .ZN(n23204) );
NAND2_X4 U33071 ( .A1(n20285), .A2(n23201), .ZN(n23202) );
NAND2_X4 U33072 ( .A1(n20247), .A2(n23202), .ZN(n23203) );
NAND2_X4 U33073 ( .A1(n23204), .A2(n23203), .ZN(n23332) );
NAND2_X4 U33074 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n23331) );
OR2_X4 U33075 ( .A1(n23332), .A2(n20209), .ZN(n23206) );
NAND2_X4 U33076 ( .A1(n20209), .A2(n23332), .ZN(n23205) );
NAND2_X4 U33077 ( .A1(n23206), .A2(n23205), .ZN(n23327) );
NAND2_X4 U33078 ( .A1(n20282), .A2(n23207), .ZN(n23212) );
NAND2_X4 U33079 ( .A1(n20318), .A2(n23208), .ZN(n23210) );
NAND2_X4 U33080 ( .A1(n23210), .A2(n23209), .ZN(n23211) );
NAND2_X4 U33081 ( .A1(n23212), .A2(n23211), .ZN(n23340) );
NAND2_X4 U33082 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n23338) );
OR2_X4 U33083 ( .A1(n23340), .A2(n20244), .ZN(n23214) );
NAND2_X4 U33084 ( .A1(n20244), .A2(n23340), .ZN(n23213) );
NAND2_X4 U33085 ( .A1(n23214), .A2(n23213), .ZN(n23324) );
NAND2_X4 U33086 ( .A1(n20319), .A2(n20355), .ZN(n23220) );
NAND2_X4 U33087 ( .A1(n23216), .A2(n23215), .ZN(n23218) );
NAND2_X4 U33088 ( .A1(n23218), .A2(n23217), .ZN(n23219) );
NAND2_X4 U33089 ( .A1(n23220), .A2(n23219), .ZN(n23348) );
NAND2_X4 U33090 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n23347) );
OR2_X4 U33091 ( .A1(n23348), .A2(n20280), .ZN(n23222) );
NAND2_X4 U33092 ( .A1(n20280), .A2(n23348), .ZN(n23221) );
NAND2_X4 U33093 ( .A1(n23222), .A2(n23221), .ZN(n23321) );
NAND2_X4 U33094 ( .A1(n20356), .A2(n23223), .ZN(n23228) );
NAND2_X4 U33095 ( .A1(n20392), .A2(n23224), .ZN(n23226) );
NAND2_X4 U33096 ( .A1(n23226), .A2(n23225), .ZN(n23227) );
NAND2_X4 U33097 ( .A1(n23228), .A2(n23227), .ZN(n23356) );
NAND2_X4 U33098 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n23354) );
OR2_X4 U33099 ( .A1(n23356), .A2(n20317), .ZN(n23230) );
NAND2_X4 U33100 ( .A1(n20317), .A2(n23356), .ZN(n23229) );
NAND2_X4 U33101 ( .A1(n23230), .A2(n23229), .ZN(n23318) );
NAND2_X4 U33102 ( .A1(n20393), .A2(n20429), .ZN(n23236) );
NAND2_X4 U33103 ( .A1(n23232), .A2(n23231), .ZN(n23234) );
NAND2_X4 U33104 ( .A1(n23234), .A2(n23233), .ZN(n23235) );
NAND2_X4 U33105 ( .A1(n23236), .A2(n23235), .ZN(n23364) );
NAND2_X4 U33106 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n23363) );
OR2_X4 U33107 ( .A1(n23364), .A2(n20354), .ZN(n23238) );
NAND2_X4 U33108 ( .A1(n20354), .A2(n23364), .ZN(n23237) );
NAND2_X4 U33109 ( .A1(n23238), .A2(n23237), .ZN(n23315) );
NAND2_X4 U33110 ( .A1(n20430), .A2(n23239), .ZN(n23244) );
NAND2_X4 U33111 ( .A1(n20467), .A2(n23240), .ZN(n23242) );
NAND2_X4 U33112 ( .A1(n23242), .A2(n23241), .ZN(n23243) );
NAND2_X4 U33113 ( .A1(n23244), .A2(n23243), .ZN(n23372) );
NAND2_X4 U33114 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n23370) );
OR2_X4 U33115 ( .A1(n23372), .A2(n20391), .ZN(n23246) );
NAND2_X4 U33116 ( .A1(n20391), .A2(n23372), .ZN(n23245) );
NAND2_X4 U33117 ( .A1(n23246), .A2(n23245), .ZN(n23312) );
NAND2_X4 U33118 ( .A1(n20468), .A2(n20505), .ZN(n23252) );
NAND2_X4 U33119 ( .A1(n23248), .A2(n23247), .ZN(n23250) );
NAND2_X4 U33120 ( .A1(n23250), .A2(n23249), .ZN(n23251) );
NAND2_X4 U33121 ( .A1(n23252), .A2(n23251), .ZN(n23380) );
NAND2_X4 U33122 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n23379) );
OR2_X4 U33123 ( .A1(n23380), .A2(n20428), .ZN(n23254) );
NAND2_X4 U33124 ( .A1(n20428), .A2(n23380), .ZN(n23253) );
NAND2_X4 U33125 ( .A1(n23254), .A2(n23253), .ZN(n23309) );
NAND2_X4 U33126 ( .A1(n20506), .A2(n23255), .ZN(n23260) );
NAND2_X4 U33127 ( .A1(n20543), .A2(n23256), .ZN(n23258) );
NAND2_X4 U33128 ( .A1(n23258), .A2(n23257), .ZN(n23259) );
NAND2_X4 U33129 ( .A1(n23260), .A2(n23259), .ZN(n23388) );
NAND2_X4 U33130 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n23386) );
OR2_X4 U33131 ( .A1(n23388), .A2(n20466), .ZN(n23262) );
NAND2_X4 U33132 ( .A1(n20466), .A2(n23388), .ZN(n23261) );
NAND2_X4 U33133 ( .A1(n23262), .A2(n23261), .ZN(n23306) );
NAND2_X4 U33134 ( .A1(n20544), .A2(n20581), .ZN(n23268) );
NAND2_X4 U33135 ( .A1(n23264), .A2(n23263), .ZN(n23266) );
NAND2_X4 U33136 ( .A1(n23266), .A2(n23265), .ZN(n23267) );
NAND2_X4 U33137 ( .A1(n23268), .A2(n23267), .ZN(n23396) );
NAND2_X4 U33138 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n23395) );
OR2_X4 U33139 ( .A1(n23396), .A2(n20504), .ZN(n23270) );
NAND2_X4 U33140 ( .A1(n20504), .A2(n23396), .ZN(n23269) );
NAND2_X4 U33141 ( .A1(n23270), .A2(n23269), .ZN(n23303) );
NAND2_X4 U33142 ( .A1(n20582), .A2(n23271), .ZN(n23276) );
NAND2_X4 U33143 ( .A1(n20618), .A2(n23272), .ZN(n23274) );
NAND2_X4 U33144 ( .A1(n23274), .A2(n23273), .ZN(n23275) );
NAND2_X4 U33145 ( .A1(n23276), .A2(n23275), .ZN(n23404) );
NAND2_X4 U33146 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n23402) );
OR2_X4 U33147 ( .A1(n23404), .A2(n20542), .ZN(n23278) );
NAND2_X4 U33148 ( .A1(n20542), .A2(n23404), .ZN(n23277) );
NAND2_X4 U33149 ( .A1(n23278), .A2(n23277), .ZN(n23300) );
NAND2_X4 U33150 ( .A1(n20619), .A2(n23279), .ZN(n23283) );
NAND2_X4 U33151 ( .A1(n20653), .A2(n23280), .ZN(n23281) );
NAND2_X4 U33152 ( .A1(n20654), .A2(n23281), .ZN(n23282) );
NAND2_X4 U33153 ( .A1(n23283), .A2(n23282), .ZN(n23412) );
NAND2_X4 U33154 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n23411) );
OR2_X4 U33155 ( .A1(n23412), .A2(n20580), .ZN(n23285) );
NAND2_X4 U33156 ( .A1(n20580), .A2(n23412), .ZN(n23284) );
NAND2_X4 U33157 ( .A1(n23285), .A2(n23284), .ZN(n23297) );
NAND2_X4 U33158 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n23419) );
NOR2_X4 U33159 ( .A1(n16200), .A2(n20771), .ZN(n23287) );
NAND2_X4 U33160 ( .A1(n23287), .A2(n23286), .ZN(n23288) );
NAND2_X4 U33161 ( .A1(n20617), .A2(n23288), .ZN(n23290) );
NAND2_X4 U33162 ( .A1(n20652), .A2(n23419), .ZN(n23289) );
NAND2_X4 U33163 ( .A1(n23290), .A2(n23289), .ZN(n23294) );
NAND2_X4 U33164 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n23291) );
NOR2_X4 U33165 ( .A1(n20771), .A2(n20675), .ZN(n23425) );
OR2_X4 U33166 ( .A1(n23291), .A2(n23425), .ZN(n23293) );
NAND2_X4 U33167 ( .A1(n23425), .A2(n23291), .ZN(n23292) );
NAND2_X4 U33168 ( .A1(n23293), .A2(n23292), .ZN(n23418) );
NAND2_X4 U33169 ( .A1(n23294), .A2(n20651), .ZN(n23296) );
OR2_X4 U33170 ( .A1(n20651), .A2(n23294), .ZN(n23295) );
NAND2_X4 U33171 ( .A1(n23296), .A2(n23295), .ZN(n23410) );
NAND2_X4 U33172 ( .A1(n23297), .A2(n20616), .ZN(n23299) );
OR2_X4 U33173 ( .A1(n20616), .A2(n23297), .ZN(n23298) );
NAND2_X4 U33174 ( .A1(n23299), .A2(n23298), .ZN(n23403) );
NAND2_X4 U33175 ( .A1(n23300), .A2(n20579), .ZN(n23302) );
OR2_X4 U33176 ( .A1(n20579), .A2(n23300), .ZN(n23301) );
NAND2_X4 U33177 ( .A1(n23302), .A2(n23301), .ZN(n23394) );
NAND2_X4 U33178 ( .A1(n23303), .A2(n20541), .ZN(n23305) );
OR2_X4 U33179 ( .A1(n20541), .A2(n23303), .ZN(n23304) );
NAND2_X4 U33180 ( .A1(n23305), .A2(n23304), .ZN(n23387) );
NAND2_X4 U33181 ( .A1(n23306), .A2(n20503), .ZN(n23308) );
OR2_X4 U33182 ( .A1(n20503), .A2(n23306), .ZN(n23307) );
NAND2_X4 U33183 ( .A1(n23308), .A2(n23307), .ZN(n23378) );
NAND2_X4 U33184 ( .A1(n23309), .A2(n20465), .ZN(n23311) );
OR2_X4 U33185 ( .A1(n20465), .A2(n23309), .ZN(n23310) );
NAND2_X4 U33186 ( .A1(n23311), .A2(n23310), .ZN(n23371) );
NAND2_X4 U33187 ( .A1(n23312), .A2(n20427), .ZN(n23314) );
OR2_X4 U33188 ( .A1(n20427), .A2(n23312), .ZN(n23313) );
NAND2_X4 U33189 ( .A1(n23314), .A2(n23313), .ZN(n23362) );
NAND2_X4 U33190 ( .A1(n23315), .A2(n20390), .ZN(n23317) );
OR2_X4 U33191 ( .A1(n20390), .A2(n23315), .ZN(n23316) );
NAND2_X4 U33192 ( .A1(n23317), .A2(n23316), .ZN(n23355) );
NAND2_X4 U33193 ( .A1(n23318), .A2(n20353), .ZN(n23320) );
OR2_X4 U33194 ( .A1(n20353), .A2(n23318), .ZN(n23319) );
NAND2_X4 U33195 ( .A1(n23320), .A2(n23319), .ZN(n23346) );
NAND2_X4 U33196 ( .A1(n23321), .A2(n20316), .ZN(n23323) );
OR2_X4 U33197 ( .A1(n20316), .A2(n23321), .ZN(n23322) );
NAND2_X4 U33198 ( .A1(n23323), .A2(n23322), .ZN(n23339) );
NAND2_X4 U33199 ( .A1(n23324), .A2(n20279), .ZN(n23326) );
OR2_X4 U33200 ( .A1(n20279), .A2(n23324), .ZN(n23325) );
NAND2_X4 U33201 ( .A1(n23326), .A2(n23325), .ZN(n23330) );
NOR2_X4 U33202 ( .A1(n23327), .A2(n20243), .ZN(n23329) );
AND2_X4 U33203 ( .A1(n20243), .A2(n23327), .ZN(n23328) );
NOR2_X4 U33204 ( .A1(n23329), .A2(n23328), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N48) );
NAND2_X4 U33205 ( .A1(n20209), .A2(n23330), .ZN(n23335) );
NAND2_X4 U33206 ( .A1(n20243), .A2(n23331), .ZN(n23333) );
NAND2_X4 U33207 ( .A1(n23333), .A2(n23332), .ZN(n23334) );
NAND2_X4 U33208 ( .A1(n23335), .A2(n23334), .ZN(n23474) );
NAND2_X4 U33209 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n23472) );
OR2_X4 U33210 ( .A1(n23474), .A2(n20171), .ZN(n23337) );
NAND2_X4 U33211 ( .A1(n20171), .A2(n23474), .ZN(n23336) );
NAND2_X4 U33212 ( .A1(n23337), .A2(n23336), .ZN(n23469) );
NAND2_X4 U33213 ( .A1(n20244), .A2(n20279), .ZN(n23343) );
NAND2_X4 U33214 ( .A1(n23339), .A2(n23338), .ZN(n23341) );
NAND2_X4 U33215 ( .A1(n23341), .A2(n23340), .ZN(n23342) );
NAND2_X4 U33216 ( .A1(n23343), .A2(n23342), .ZN(n23482) );
NAND2_X4 U33217 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n23481) );
OR2_X4 U33218 ( .A1(n23482), .A2(n20206), .ZN(n23345) );
NAND2_X4 U33219 ( .A1(n20206), .A2(n23482), .ZN(n23344) );
NAND2_X4 U33220 ( .A1(n23345), .A2(n23344), .ZN(n23466) );
NAND2_X4 U33221 ( .A1(n20280), .A2(n23346), .ZN(n23351) );
NAND2_X4 U33222 ( .A1(n20316), .A2(n23347), .ZN(n23349) );
NAND2_X4 U33223 ( .A1(n23349), .A2(n23348), .ZN(n23350) );
NAND2_X4 U33224 ( .A1(n23351), .A2(n23350), .ZN(n23490) );
NAND2_X4 U33225 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n23488) );
OR2_X4 U33226 ( .A1(n23490), .A2(n20242), .ZN(n23353) );
NAND2_X4 U33227 ( .A1(n20242), .A2(n23490), .ZN(n23352) );
NAND2_X4 U33228 ( .A1(n23353), .A2(n23352), .ZN(n23463) );
NAND2_X4 U33229 ( .A1(n20317), .A2(n20353), .ZN(n23359) );
NAND2_X4 U33230 ( .A1(n23355), .A2(n23354), .ZN(n23357) );
NAND2_X4 U33231 ( .A1(n23357), .A2(n23356), .ZN(n23358) );
NAND2_X4 U33232 ( .A1(n23359), .A2(n23358), .ZN(n23498) );
NAND2_X4 U33233 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n23497) );
OR2_X4 U33234 ( .A1(n23498), .A2(n20278), .ZN(n23361) );
NAND2_X4 U33235 ( .A1(n20278), .A2(n23498), .ZN(n23360) );
NAND2_X4 U33236 ( .A1(n23361), .A2(n23360), .ZN(n23460) );
NAND2_X4 U33237 ( .A1(n20354), .A2(n23362), .ZN(n23367) );
NAND2_X4 U33238 ( .A1(n20390), .A2(n23363), .ZN(n23365) );
NAND2_X4 U33239 ( .A1(n23365), .A2(n23364), .ZN(n23366) );
NAND2_X4 U33240 ( .A1(n23367), .A2(n23366), .ZN(n23506) );
NAND2_X4 U33241 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n23504) );
OR2_X4 U33242 ( .A1(n23506), .A2(n20315), .ZN(n23369) );
NAND2_X4 U33243 ( .A1(n20315), .A2(n23506), .ZN(n23368) );
NAND2_X4 U33244 ( .A1(n23369), .A2(n23368), .ZN(n23457) );
NAND2_X4 U33245 ( .A1(n20391), .A2(n20427), .ZN(n23375) );
NAND2_X4 U33246 ( .A1(n23371), .A2(n23370), .ZN(n23373) );
NAND2_X4 U33247 ( .A1(n23373), .A2(n23372), .ZN(n23374) );
NAND2_X4 U33248 ( .A1(n23375), .A2(n23374), .ZN(n23514) );
NAND2_X4 U33249 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n23513) );
OR2_X4 U33250 ( .A1(n23514), .A2(n20352), .ZN(n23377) );
NAND2_X4 U33251 ( .A1(n20352), .A2(n23514), .ZN(n23376) );
NAND2_X4 U33252 ( .A1(n23377), .A2(n23376), .ZN(n23454) );
NAND2_X4 U33253 ( .A1(n20428), .A2(n23378), .ZN(n23383) );
NAND2_X4 U33254 ( .A1(n20465), .A2(n23379), .ZN(n23381) );
NAND2_X4 U33255 ( .A1(n23381), .A2(n23380), .ZN(n23382) );
NAND2_X4 U33256 ( .A1(n23383), .A2(n23382), .ZN(n23522) );
NAND2_X4 U33257 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n23520) );
OR2_X4 U33258 ( .A1(n23522), .A2(n20389), .ZN(n23385) );
NAND2_X4 U33259 ( .A1(n20389), .A2(n23522), .ZN(n23384) );
NAND2_X4 U33260 ( .A1(n23385), .A2(n23384), .ZN(n23451) );
NAND2_X4 U33261 ( .A1(n20466), .A2(n20503), .ZN(n23391) );
NAND2_X4 U33262 ( .A1(n23387), .A2(n23386), .ZN(n23389) );
NAND2_X4 U33263 ( .A1(n23389), .A2(n23388), .ZN(n23390) );
NAND2_X4 U33264 ( .A1(n23391), .A2(n23390), .ZN(n23530) );
NAND2_X4 U33265 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n23529) );
OR2_X4 U33266 ( .A1(n23530), .A2(n20426), .ZN(n23393) );
NAND2_X4 U33267 ( .A1(n20426), .A2(n23530), .ZN(n23392) );
NAND2_X4 U33268 ( .A1(n23393), .A2(n23392), .ZN(n23448) );
NAND2_X4 U33269 ( .A1(n20504), .A2(n23394), .ZN(n23399) );
NAND2_X4 U33270 ( .A1(n20541), .A2(n23395), .ZN(n23397) );
NAND2_X4 U33271 ( .A1(n23397), .A2(n23396), .ZN(n23398) );
NAND2_X4 U33272 ( .A1(n23399), .A2(n23398), .ZN(n23538) );
NAND2_X4 U33273 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n23536) );
OR2_X4 U33274 ( .A1(n23538), .A2(n20464), .ZN(n23401) );
NAND2_X4 U33275 ( .A1(n20464), .A2(n23538), .ZN(n23400) );
NAND2_X4 U33276 ( .A1(n23401), .A2(n23400), .ZN(n23445) );
NAND2_X4 U33277 ( .A1(n20542), .A2(n20579), .ZN(n23407) );
NAND2_X4 U33278 ( .A1(n23403), .A2(n23402), .ZN(n23405) );
NAND2_X4 U33279 ( .A1(n23405), .A2(n23404), .ZN(n23406) );
NAND2_X4 U33280 ( .A1(n23407), .A2(n23406), .ZN(n23546) );
NAND2_X4 U33281 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n23545) );
OR2_X4 U33282 ( .A1(n23546), .A2(n20502), .ZN(n23409) );
NAND2_X4 U33283 ( .A1(n20502), .A2(n23546), .ZN(n23408) );
NAND2_X4 U33284 ( .A1(n23409), .A2(n23408), .ZN(n23442) );
NAND2_X4 U33285 ( .A1(n20580), .A2(n23410), .ZN(n23415) );
NAND2_X4 U33286 ( .A1(n20616), .A2(n23411), .ZN(n23413) );
NAND2_X4 U33287 ( .A1(n23413), .A2(n23412), .ZN(n23414) );
NAND2_X4 U33288 ( .A1(n23415), .A2(n23414), .ZN(n23554) );
NAND2_X4 U33289 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n23552) );
OR2_X4 U33290 ( .A1(n23554), .A2(n20540), .ZN(n23417) );
NAND2_X4 U33291 ( .A1(n20540), .A2(n23554), .ZN(n23416) );
NAND2_X4 U33292 ( .A1(n23417), .A2(n23416), .ZN(n23439) );
NAND2_X4 U33293 ( .A1(n20617), .A2(n23418), .ZN(n23422) );
NAND2_X4 U33294 ( .A1(n20651), .A2(n23419), .ZN(n23420) );
NAND2_X4 U33295 ( .A1(n20652), .A2(n23420), .ZN(n23421) );
NAND2_X4 U33296 ( .A1(n23422), .A2(n23421), .ZN(n23562) );
NAND2_X4 U33297 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n23561) );
OR2_X4 U33298 ( .A1(n23562), .A2(n20578), .ZN(n23424) );
NAND2_X4 U33299 ( .A1(n20578), .A2(n23562), .ZN(n23423) );
NAND2_X4 U33300 ( .A1(n23424), .A2(n23423), .ZN(n23436) );
NAND2_X4 U33301 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n23569) );
NOR2_X4 U33302 ( .A1(n16200), .A2(n20768), .ZN(n23426) );
NAND2_X4 U33303 ( .A1(n23426), .A2(n23425), .ZN(n23427) );
NAND2_X4 U33304 ( .A1(n20615), .A2(n23427), .ZN(n23429) );
NAND2_X4 U33305 ( .A1(n20650), .A2(n23569), .ZN(n23428) );
NAND2_X4 U33306 ( .A1(n23429), .A2(n23428), .ZN(n23433) );
NAND2_X4 U33307 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n23430) );
NOR2_X4 U33308 ( .A1(n20768), .A2(n20675), .ZN(n23575) );
OR2_X4 U33309 ( .A1(n23430), .A2(n23575), .ZN(n23432) );
NAND2_X4 U33310 ( .A1(n23575), .A2(n23430), .ZN(n23431) );
NAND2_X4 U33311 ( .A1(n23432), .A2(n23431), .ZN(n23568) );
NAND2_X4 U33312 ( .A1(n23433), .A2(n20649), .ZN(n23435) );
OR2_X4 U33313 ( .A1(n20649), .A2(n23433), .ZN(n23434) );
NAND2_X4 U33314 ( .A1(n23435), .A2(n23434), .ZN(n23560) );
NAND2_X4 U33315 ( .A1(n23436), .A2(n20614), .ZN(n23438) );
OR2_X4 U33316 ( .A1(n20614), .A2(n23436), .ZN(n23437) );
NAND2_X4 U33317 ( .A1(n23438), .A2(n23437), .ZN(n23553) );
NAND2_X4 U33318 ( .A1(n23439), .A2(n20577), .ZN(n23441) );
OR2_X4 U33319 ( .A1(n20577), .A2(n23439), .ZN(n23440) );
NAND2_X4 U33320 ( .A1(n23441), .A2(n23440), .ZN(n23544) );
NAND2_X4 U33321 ( .A1(n23442), .A2(n20539), .ZN(n23444) );
OR2_X4 U33322 ( .A1(n20539), .A2(n23442), .ZN(n23443) );
NAND2_X4 U33323 ( .A1(n23444), .A2(n23443), .ZN(n23537) );
NAND2_X4 U33324 ( .A1(n23445), .A2(n20501), .ZN(n23447) );
OR2_X4 U33325 ( .A1(n20501), .A2(n23445), .ZN(n23446) );
NAND2_X4 U33326 ( .A1(n23447), .A2(n23446), .ZN(n23528) );
NAND2_X4 U33327 ( .A1(n23448), .A2(n20463), .ZN(n23450) );
OR2_X4 U33328 ( .A1(n20463), .A2(n23448), .ZN(n23449) );
NAND2_X4 U33329 ( .A1(n23450), .A2(n23449), .ZN(n23521) );
NAND2_X4 U33330 ( .A1(n23451), .A2(n20425), .ZN(n23453) );
OR2_X4 U33331 ( .A1(n20425), .A2(n23451), .ZN(n23452) );
NAND2_X4 U33332 ( .A1(n23453), .A2(n23452), .ZN(n23512) );
NAND2_X4 U33333 ( .A1(n23454), .A2(n20388), .ZN(n23456) );
OR2_X4 U33334 ( .A1(n20388), .A2(n23454), .ZN(n23455) );
NAND2_X4 U33335 ( .A1(n23456), .A2(n23455), .ZN(n23505) );
NAND2_X4 U33336 ( .A1(n23457), .A2(n20351), .ZN(n23459) );
OR2_X4 U33337 ( .A1(n20351), .A2(n23457), .ZN(n23458) );
NAND2_X4 U33338 ( .A1(n23459), .A2(n23458), .ZN(n23496) );
NAND2_X4 U33339 ( .A1(n23460), .A2(n20314), .ZN(n23462) );
OR2_X4 U33340 ( .A1(n20314), .A2(n23460), .ZN(n23461) );
NAND2_X4 U33341 ( .A1(n23462), .A2(n23461), .ZN(n23489) );
NAND2_X4 U33342 ( .A1(n23463), .A2(n20277), .ZN(n23465) );
OR2_X4 U33343 ( .A1(n20277), .A2(n23463), .ZN(n23464) );
NAND2_X4 U33344 ( .A1(n23465), .A2(n23464), .ZN(n23480) );
NAND2_X4 U33345 ( .A1(n23466), .A2(n16331), .ZN(n23468) );
OR2_X4 U33346 ( .A1(n16331), .A2(n23466), .ZN(n23467) );
NAND2_X4 U33347 ( .A1(n23468), .A2(n23467), .ZN(n23473) );
NAND2_X4 U33348 ( .A1(n23469), .A2(n20205), .ZN(n23471) );
OR2_X4 U33349 ( .A1(n20205), .A2(n23469), .ZN(n23470) );
NAND2_X4 U33350 ( .A1(n23471), .A2(n23470), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N49) );
NAND2_X4 U33351 ( .A1(n20171), .A2(n20205), .ZN(n23477) );
NAND2_X4 U33352 ( .A1(n23473), .A2(n23472), .ZN(n23475) );
NAND2_X4 U33353 ( .A1(n23475), .A2(n23474), .ZN(n23476) );
NAND2_X4 U33354 ( .A1(n23477), .A2(n23476), .ZN(n23781) );
NAND2_X4 U33355 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n23780) );
OR2_X4 U33356 ( .A1(n23781), .A2(n20109), .ZN(n23479) );
NAND2_X4 U33357 ( .A1(n20109), .A2(n23781), .ZN(n23478) );
NAND2_X4 U33358 ( .A1(n23479), .A2(n23478), .ZN(n23622) );
NAND2_X4 U33359 ( .A1(n20206), .A2(n23480), .ZN(n23485) );
NAND2_X4 U33360 ( .A1(n20241), .A2(n23481), .ZN(n23483) );
NAND2_X4 U33361 ( .A1(n23483), .A2(n23482), .ZN(n23484) );
NAND2_X4 U33362 ( .A1(n23485), .A2(n23484), .ZN(n23629) );
NAND2_X4 U33363 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n23627) );
OR2_X4 U33364 ( .A1(n23629), .A2(n20168), .ZN(n23487) );
NAND2_X4 U33365 ( .A1(n20168), .A2(n23629), .ZN(n23486) );
NAND2_X4 U33366 ( .A1(n23487), .A2(n23486), .ZN(n23619) );
NAND2_X4 U33367 ( .A1(n20242), .A2(n20277), .ZN(n23493) );
NAND2_X4 U33368 ( .A1(n23489), .A2(n23488), .ZN(n23491) );
NAND2_X4 U33369 ( .A1(n23491), .A2(n23490), .ZN(n23492) );
NAND2_X4 U33370 ( .A1(n23493), .A2(n23492), .ZN(n23637) );
NAND2_X4 U33371 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n23636) );
OR2_X4 U33372 ( .A1(n23637), .A2(n20204), .ZN(n23495) );
NAND2_X4 U33373 ( .A1(n20204), .A2(n23637), .ZN(n23494) );
NAND2_X4 U33374 ( .A1(n23495), .A2(n23494), .ZN(n23616) );
NAND2_X4 U33375 ( .A1(n20278), .A2(n23496), .ZN(n23501) );
NAND2_X4 U33376 ( .A1(n16198), .A2(n23497), .ZN(n23499) );
NAND2_X4 U33377 ( .A1(n23499), .A2(n23498), .ZN(n23500) );
NAND2_X4 U33378 ( .A1(n23501), .A2(n23500), .ZN(n23645) );
NAND2_X4 U33379 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n23643) );
OR2_X4 U33380 ( .A1(n23645), .A2(n20240), .ZN(n23503) );
NAND2_X4 U33381 ( .A1(n20240), .A2(n23645), .ZN(n23502) );
NAND2_X4 U33382 ( .A1(n23503), .A2(n23502), .ZN(n23613) );
NAND2_X4 U33383 ( .A1(n20315), .A2(n20351), .ZN(n23509) );
NAND2_X4 U33384 ( .A1(n23505), .A2(n23504), .ZN(n23507) );
NAND2_X4 U33385 ( .A1(n23507), .A2(n23506), .ZN(n23508) );
NAND2_X4 U33386 ( .A1(n23509), .A2(n23508), .ZN(n23653) );
NAND2_X4 U33387 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n23652) );
OR2_X4 U33388 ( .A1(n23653), .A2(n20276), .ZN(n23511) );
NAND2_X4 U33389 ( .A1(n20276), .A2(n23653), .ZN(n23510) );
NAND2_X4 U33390 ( .A1(n23511), .A2(n23510), .ZN(n23610) );
NAND2_X4 U33391 ( .A1(n20352), .A2(n23512), .ZN(n23517) );
NAND2_X4 U33392 ( .A1(n20388), .A2(n23513), .ZN(n23515) );
NAND2_X4 U33393 ( .A1(n23515), .A2(n23514), .ZN(n23516) );
NAND2_X4 U33394 ( .A1(n23517), .A2(n23516), .ZN(n23661) );
NAND2_X4 U33395 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n23659) );
OR2_X4 U33396 ( .A1(n23661), .A2(n20313), .ZN(n23519) );
NAND2_X4 U33397 ( .A1(n20313), .A2(n23661), .ZN(n23518) );
NAND2_X4 U33398 ( .A1(n23519), .A2(n23518), .ZN(n23607) );
NAND2_X4 U33399 ( .A1(n20389), .A2(n20425), .ZN(n23525) );
NAND2_X4 U33400 ( .A1(n23521), .A2(n23520), .ZN(n23523) );
NAND2_X4 U33401 ( .A1(n23523), .A2(n23522), .ZN(n23524) );
NAND2_X4 U33402 ( .A1(n23525), .A2(n23524), .ZN(n23669) );
NAND2_X4 U33403 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n23668) );
OR2_X4 U33404 ( .A1(n23669), .A2(n20350), .ZN(n23527) );
NAND2_X4 U33405 ( .A1(n20350), .A2(n23669), .ZN(n23526) );
NAND2_X4 U33406 ( .A1(n23527), .A2(n23526), .ZN(n23604) );
NAND2_X4 U33407 ( .A1(n20426), .A2(n23528), .ZN(n23533) );
NAND2_X4 U33408 ( .A1(n20463), .A2(n23529), .ZN(n23531) );
NAND2_X4 U33409 ( .A1(n23531), .A2(n23530), .ZN(n23532) );
NAND2_X4 U33410 ( .A1(n23533), .A2(n23532), .ZN(n23677) );
NAND2_X4 U33411 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n23675) );
OR2_X4 U33412 ( .A1(n23677), .A2(n20387), .ZN(n23535) );
NAND2_X4 U33413 ( .A1(n20387), .A2(n23677), .ZN(n23534) );
NAND2_X4 U33414 ( .A1(n23535), .A2(n23534), .ZN(n23601) );
NAND2_X4 U33415 ( .A1(n20464), .A2(n20501), .ZN(n23541) );
NAND2_X4 U33416 ( .A1(n23537), .A2(n23536), .ZN(n23539) );
NAND2_X4 U33417 ( .A1(n23539), .A2(n23538), .ZN(n23540) );
NAND2_X4 U33418 ( .A1(n23541), .A2(n23540), .ZN(n23685) );
NAND2_X4 U33419 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n23684) );
OR2_X4 U33420 ( .A1(n23685), .A2(n20424), .ZN(n23543) );
NAND2_X4 U33421 ( .A1(n20424), .A2(n23685), .ZN(n23542) );
NAND2_X4 U33422 ( .A1(n23543), .A2(n23542), .ZN(n23598) );
NAND2_X4 U33423 ( .A1(n20502), .A2(n23544), .ZN(n23549) );
NAND2_X4 U33424 ( .A1(n20539), .A2(n23545), .ZN(n23547) );
NAND2_X4 U33425 ( .A1(n23547), .A2(n23546), .ZN(n23548) );
NAND2_X4 U33426 ( .A1(n23549), .A2(n23548), .ZN(n23693) );
NAND2_X4 U33427 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n23691) );
OR2_X4 U33428 ( .A1(n23693), .A2(n20462), .ZN(n23551) );
NAND2_X4 U33429 ( .A1(n20462), .A2(n23693), .ZN(n23550) );
NAND2_X4 U33430 ( .A1(n23551), .A2(n23550), .ZN(n23595) );
NAND2_X4 U33431 ( .A1(n20540), .A2(n20577), .ZN(n23557) );
NAND2_X4 U33432 ( .A1(n23553), .A2(n23552), .ZN(n23555) );
NAND2_X4 U33433 ( .A1(n23555), .A2(n23554), .ZN(n23556) );
NAND2_X4 U33434 ( .A1(n23557), .A2(n23556), .ZN(n23701) );
NAND2_X4 U33435 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n23700) );
OR2_X4 U33436 ( .A1(n23701), .A2(n20500), .ZN(n23559) );
NAND2_X4 U33437 ( .A1(n20500), .A2(n23701), .ZN(n23558) );
NAND2_X4 U33438 ( .A1(n23559), .A2(n23558), .ZN(n23592) );
NAND2_X4 U33439 ( .A1(n20578), .A2(n23560), .ZN(n23565) );
NAND2_X4 U33440 ( .A1(n20614), .A2(n23561), .ZN(n23563) );
NAND2_X4 U33441 ( .A1(n23563), .A2(n23562), .ZN(n23564) );
NAND2_X4 U33442 ( .A1(n23565), .A2(n23564), .ZN(n23709) );
NAND2_X4 U33443 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n23707) );
OR2_X4 U33444 ( .A1(n23709), .A2(n20538), .ZN(n23567) );
NAND2_X4 U33445 ( .A1(n20538), .A2(n23709), .ZN(n23566) );
NAND2_X4 U33446 ( .A1(n23567), .A2(n23566), .ZN(n23589) );
NAND2_X4 U33447 ( .A1(n20615), .A2(n23568), .ZN(n23572) );
NAND2_X4 U33448 ( .A1(n20649), .A2(n23569), .ZN(n23570) );
NAND2_X4 U33449 ( .A1(n20650), .A2(n23570), .ZN(n23571) );
NAND2_X4 U33450 ( .A1(n23572), .A2(n23571), .ZN(n23717) );
NAND2_X4 U33451 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n23716) );
OR2_X4 U33452 ( .A1(n23717), .A2(n20576), .ZN(n23574) );
NAND2_X4 U33453 ( .A1(n20576), .A2(n23717), .ZN(n23573) );
NAND2_X4 U33454 ( .A1(n23574), .A2(n23573), .ZN(n23586) );
NAND2_X4 U33455 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n23724) );
NOR2_X4 U33456 ( .A1(n16200), .A2(n20765), .ZN(n23576) );
NAND2_X4 U33457 ( .A1(n23576), .A2(n23575), .ZN(n23577) );
NAND2_X4 U33458 ( .A1(n20613), .A2(n23577), .ZN(n23579) );
NAND2_X4 U33459 ( .A1(n20648), .A2(n23724), .ZN(n23578) );
NAND2_X4 U33460 ( .A1(n23579), .A2(n23578), .ZN(n23583) );
NAND2_X4 U33461 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n23580) );
NOR2_X4 U33462 ( .A1(n20765), .A2(n20675), .ZN(n23730) );
OR2_X4 U33463 ( .A1(n23580), .A2(n23730), .ZN(n23582) );
NAND2_X4 U33464 ( .A1(n23730), .A2(n23580), .ZN(n23581) );
NAND2_X4 U33465 ( .A1(n23582), .A2(n23581), .ZN(n23723) );
NAND2_X4 U33466 ( .A1(n23583), .A2(n20647), .ZN(n23585) );
OR2_X4 U33467 ( .A1(n20647), .A2(n23583), .ZN(n23584) );
NAND2_X4 U33468 ( .A1(n23585), .A2(n23584), .ZN(n23715) );
NAND2_X4 U33469 ( .A1(n23586), .A2(n20612), .ZN(n23588) );
OR2_X4 U33470 ( .A1(n20612), .A2(n23586), .ZN(n23587) );
NAND2_X4 U33471 ( .A1(n23588), .A2(n23587), .ZN(n23708) );
NAND2_X4 U33472 ( .A1(n23589), .A2(n20575), .ZN(n23591) );
OR2_X4 U33473 ( .A1(n20575), .A2(n23589), .ZN(n23590) );
NAND2_X4 U33474 ( .A1(n23591), .A2(n23590), .ZN(n23699) );
NAND2_X4 U33475 ( .A1(n23592), .A2(n20537), .ZN(n23594) );
OR2_X4 U33476 ( .A1(n20537), .A2(n23592), .ZN(n23593) );
NAND2_X4 U33477 ( .A1(n23594), .A2(n23593), .ZN(n23692) );
NAND2_X4 U33478 ( .A1(n23595), .A2(n20499), .ZN(n23597) );
OR2_X4 U33479 ( .A1(n20499), .A2(n23595), .ZN(n23596) );
NAND2_X4 U33480 ( .A1(n23597), .A2(n23596), .ZN(n23683) );
NAND2_X4 U33481 ( .A1(n23598), .A2(n20461), .ZN(n23600) );
OR2_X4 U33482 ( .A1(n20461), .A2(n23598), .ZN(n23599) );
NAND2_X4 U33483 ( .A1(n23600), .A2(n23599), .ZN(n23676) );
NAND2_X4 U33484 ( .A1(n23601), .A2(n20423), .ZN(n23603) );
OR2_X4 U33485 ( .A1(n20423), .A2(n23601), .ZN(n23602) );
NAND2_X4 U33486 ( .A1(n23603), .A2(n23602), .ZN(n23667) );
NAND2_X4 U33487 ( .A1(n23604), .A2(n20386), .ZN(n23606) );
OR2_X4 U33488 ( .A1(n20386), .A2(n23604), .ZN(n23605) );
NAND2_X4 U33489 ( .A1(n23606), .A2(n23605), .ZN(n23660) );
NAND2_X4 U33490 ( .A1(n23607), .A2(n20349), .ZN(n23609) );
OR2_X4 U33491 ( .A1(n20349), .A2(n23607), .ZN(n23608) );
NAND2_X4 U33492 ( .A1(n23609), .A2(n23608), .ZN(n23651) );
NAND2_X4 U33493 ( .A1(n23610), .A2(n20312), .ZN(n23612) );
OR2_X4 U33494 ( .A1(n20312), .A2(n23610), .ZN(n23611) );
NAND2_X4 U33495 ( .A1(n23612), .A2(n23611), .ZN(n23644) );
NAND2_X4 U33496 ( .A1(n23613), .A2(n20275), .ZN(n23615) );
OR2_X4 U33497 ( .A1(n20275), .A2(n23613), .ZN(n23614) );
NAND2_X4 U33498 ( .A1(n23615), .A2(n23614), .ZN(n23635) );
NAND2_X4 U33499 ( .A1(n23616), .A2(n20239), .ZN(n23618) );
OR2_X4 U33500 ( .A1(n20239), .A2(n23616), .ZN(n23617) );
NAND2_X4 U33501 ( .A1(n23618), .A2(n23617), .ZN(n23628) );
NAND2_X4 U33502 ( .A1(n23619), .A2(n20203), .ZN(n23621) );
OR2_X4 U33503 ( .A1(n20203), .A2(n23619), .ZN(n23620) );
NAND2_X4 U33504 ( .A1(n23621), .A2(n23620), .ZN(n23779) );
NOR2_X4 U33505 ( .A1(n23622), .A2(n20167), .ZN(n23624) );
AND2_X4 U33506 ( .A1(n20167), .A2(n23622), .ZN(n23623) );
NOR2_X4 U33507 ( .A1(n23624), .A2(n23623), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N50) );
NAND2_X4 U33508 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_sign_a), .A2(n20762), .ZN(n23626) );
NAND2_X4 U33509 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_sign_b), .A2(n20084), .ZN(n23625) );
NAND2_X4 U33510 ( .A1(n23626), .A2(n23625), .ZN(n25191) );
NAND2_X4 U33511 ( .A1(n20168), .A2(n20203), .ZN(n23632) );
NAND2_X4 U33512 ( .A1(n23628), .A2(n23627), .ZN(n23630) );
NAND2_X4 U33513 ( .A1(n23630), .A2(n23629), .ZN(n23631) );
NAND2_X4 U33514 ( .A1(n23632), .A2(n23631), .ZN(n23941) );
NAND2_X4 U33515 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n23940) );
OR2_X4 U33516 ( .A1(n23941), .A2(n20106), .ZN(n23634) );
NAND2_X4 U33517 ( .A1(n20106), .A2(n23941), .ZN(n23633) );
NAND2_X4 U33518 ( .A1(n23634), .A2(n23633), .ZN(n23776) );
NAND2_X4 U33519 ( .A1(n20204), .A2(n23635), .ZN(n23640) );
NAND2_X4 U33520 ( .A1(n16199), .A2(n23636), .ZN(n23638) );
NAND2_X4 U33521 ( .A1(n23638), .A2(n23637), .ZN(n23639) );
NAND2_X4 U33522 ( .A1(n23640), .A2(n23639), .ZN(n23793) );
NAND2_X4 U33523 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n23791) );
OR2_X4 U33524 ( .A1(n23793), .A2(n20166), .ZN(n23642) );
NAND2_X4 U33525 ( .A1(n20166), .A2(n23793), .ZN(n23641) );
NAND2_X4 U33526 ( .A1(n23642), .A2(n23641), .ZN(n23773) );
NAND2_X4 U33527 ( .A1(n20240), .A2(n20275), .ZN(n23648) );
NAND2_X4 U33528 ( .A1(n23644), .A2(n23643), .ZN(n23646) );
NAND2_X4 U33529 ( .A1(n23646), .A2(n23645), .ZN(n23647) );
NAND2_X4 U33530 ( .A1(n23648), .A2(n23647), .ZN(n23801) );
NAND2_X4 U33531 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n23800) );
OR2_X4 U33532 ( .A1(n23801), .A2(n20202), .ZN(n23650) );
NAND2_X4 U33533 ( .A1(n20202), .A2(n23801), .ZN(n23649) );
NAND2_X4 U33534 ( .A1(n23650), .A2(n23649), .ZN(n23770) );
NAND2_X4 U33535 ( .A1(n20276), .A2(n23651), .ZN(n23656) );
NAND2_X4 U33536 ( .A1(n20312), .A2(n23652), .ZN(n23654) );
NAND2_X4 U33537 ( .A1(n23654), .A2(n23653), .ZN(n23655) );
NAND2_X4 U33538 ( .A1(n23656), .A2(n23655), .ZN(n23809) );
NAND2_X4 U33539 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n23807) );
OR2_X4 U33540 ( .A1(n23809), .A2(n20238), .ZN(n23658) );
NAND2_X4 U33541 ( .A1(n20238), .A2(n23809), .ZN(n23657) );
NAND2_X4 U33542 ( .A1(n23658), .A2(n23657), .ZN(n23767) );
NAND2_X4 U33543 ( .A1(n20313), .A2(n20349), .ZN(n23664) );
NAND2_X4 U33544 ( .A1(n23660), .A2(n23659), .ZN(n23662) );
NAND2_X4 U33545 ( .A1(n23662), .A2(n23661), .ZN(n23663) );
NAND2_X4 U33546 ( .A1(n23664), .A2(n23663), .ZN(n23817) );
NAND2_X4 U33547 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n23816) );
OR2_X4 U33548 ( .A1(n23817), .A2(n20274), .ZN(n23666) );
NAND2_X4 U33549 ( .A1(n20274), .A2(n23817), .ZN(n23665) );
NAND2_X4 U33550 ( .A1(n23666), .A2(n23665), .ZN(n23764) );
NAND2_X4 U33551 ( .A1(n20350), .A2(n23667), .ZN(n23672) );
NAND2_X4 U33552 ( .A1(n20386), .A2(n23668), .ZN(n23670) );
NAND2_X4 U33553 ( .A1(n23670), .A2(n23669), .ZN(n23671) );
NAND2_X4 U33554 ( .A1(n23672), .A2(n23671), .ZN(n23825) );
NAND2_X4 U33555 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n23823) );
OR2_X4 U33556 ( .A1(n23825), .A2(n20311), .ZN(n23674) );
NAND2_X4 U33557 ( .A1(n20311), .A2(n23825), .ZN(n23673) );
NAND2_X4 U33558 ( .A1(n23674), .A2(n23673), .ZN(n23761) );
NAND2_X4 U33559 ( .A1(n20387), .A2(n20423), .ZN(n23680) );
NAND2_X4 U33560 ( .A1(n23676), .A2(n23675), .ZN(n23678) );
NAND2_X4 U33561 ( .A1(n23678), .A2(n23677), .ZN(n23679) );
NAND2_X4 U33562 ( .A1(n23680), .A2(n23679), .ZN(n23833) );
NAND2_X4 U33563 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n23832) );
OR2_X4 U33564 ( .A1(n23833), .A2(n20348), .ZN(n23682) );
NAND2_X4 U33565 ( .A1(n20348), .A2(n23833), .ZN(n23681) );
NAND2_X4 U33566 ( .A1(n23682), .A2(n23681), .ZN(n23758) );
NAND2_X4 U33567 ( .A1(n20424), .A2(n23683), .ZN(n23688) );
NAND2_X4 U33568 ( .A1(n20461), .A2(n23684), .ZN(n23686) );
NAND2_X4 U33569 ( .A1(n23686), .A2(n23685), .ZN(n23687) );
NAND2_X4 U33570 ( .A1(n23688), .A2(n23687), .ZN(n23841) );
NAND2_X4 U33571 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n23839) );
OR2_X4 U33572 ( .A1(n23841), .A2(n20385), .ZN(n23690) );
NAND2_X4 U33573 ( .A1(n20385), .A2(n23841), .ZN(n23689) );
NAND2_X4 U33574 ( .A1(n23690), .A2(n23689), .ZN(n23755) );
NAND2_X4 U33575 ( .A1(n20462), .A2(n20499), .ZN(n23696) );
NAND2_X4 U33576 ( .A1(n23692), .A2(n23691), .ZN(n23694) );
NAND2_X4 U33577 ( .A1(n23694), .A2(n23693), .ZN(n23695) );
NAND2_X4 U33578 ( .A1(n23696), .A2(n23695), .ZN(n23849) );
NAND2_X4 U33579 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n23848) );
OR2_X4 U33580 ( .A1(n23849), .A2(n20422), .ZN(n23698) );
NAND2_X4 U33581 ( .A1(n20422), .A2(n23849), .ZN(n23697) );
NAND2_X4 U33582 ( .A1(n23698), .A2(n23697), .ZN(n23752) );
NAND2_X4 U33583 ( .A1(n20500), .A2(n23699), .ZN(n23704) );
NAND2_X4 U33584 ( .A1(n20537), .A2(n23700), .ZN(n23702) );
NAND2_X4 U33585 ( .A1(n23702), .A2(n23701), .ZN(n23703) );
NAND2_X4 U33586 ( .A1(n23704), .A2(n23703), .ZN(n23857) );
NAND2_X4 U33587 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n23855) );
OR2_X4 U33588 ( .A1(n23857), .A2(n20460), .ZN(n23706) );
NAND2_X4 U33589 ( .A1(n20460), .A2(n23857), .ZN(n23705) );
NAND2_X4 U33590 ( .A1(n23706), .A2(n23705), .ZN(n23749) );
NAND2_X4 U33591 ( .A1(n20538), .A2(n20575), .ZN(n23712) );
NAND2_X4 U33592 ( .A1(n23708), .A2(n23707), .ZN(n23710) );
NAND2_X4 U33593 ( .A1(n23710), .A2(n23709), .ZN(n23711) );
NAND2_X4 U33594 ( .A1(n23712), .A2(n23711), .ZN(n23865) );
NAND2_X4 U33595 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n23864) );
OR2_X4 U33596 ( .A1(n23865), .A2(n20498), .ZN(n23714) );
NAND2_X4 U33597 ( .A1(n20498), .A2(n23865), .ZN(n23713) );
NAND2_X4 U33598 ( .A1(n23714), .A2(n23713), .ZN(n23746) );
NAND2_X4 U33599 ( .A1(n20576), .A2(n23715), .ZN(n23720) );
NAND2_X4 U33600 ( .A1(n20612), .A2(n23716), .ZN(n23718) );
NAND2_X4 U33601 ( .A1(n23718), .A2(n23717), .ZN(n23719) );
NAND2_X4 U33602 ( .A1(n23720), .A2(n23719), .ZN(n23873) );
NAND2_X4 U33603 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n23871) );
OR2_X4 U33604 ( .A1(n23873), .A2(n20536), .ZN(n23722) );
NAND2_X4 U33605 ( .A1(n20536), .A2(n23873), .ZN(n23721) );
NAND2_X4 U33606 ( .A1(n23722), .A2(n23721), .ZN(n23743) );
NAND2_X4 U33607 ( .A1(n20613), .A2(n23723), .ZN(n23727) );
NAND2_X4 U33608 ( .A1(n20647), .A2(n23724), .ZN(n23725) );
NAND2_X4 U33609 ( .A1(n20648), .A2(n23725), .ZN(n23726) );
NAND2_X4 U33610 ( .A1(n23727), .A2(n23726), .ZN(n23881) );
NAND2_X4 U33611 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n23880) );
OR2_X4 U33612 ( .A1(n23881), .A2(n20574), .ZN(n23729) );
NAND2_X4 U33613 ( .A1(n20574), .A2(n23881), .ZN(n23728) );
NAND2_X4 U33614 ( .A1(n23729), .A2(n23728), .ZN(n23740) );
AND2_X4 U33615 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n23888) );
AND2_X4 U33616 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .A2(n23730), .ZN(n23731) );
NAND2_X4 U33617 ( .A1(n23731), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n23889) );
NAND2_X4 U33618 ( .A1(n23888), .A2(n23889), .ZN(n23733) );
OR2_X4 U33619 ( .A1(n23889), .A2(n23888), .ZN(n23732) );
AND2_X4 U33620 ( .A1(n23733), .A2(n23732), .ZN(n23737) );
NOR2_X4 U33621 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n23734) );
NAND2_X4 U33622 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_1), .ZN(n23893) );
NAND2_X4 U33623 ( .A1(n23734), .A2(n23893), .ZN(n23736) );
OR2_X4 U33624 ( .A1(n23893), .A2(n23734), .ZN(n23735) );
NAND2_X4 U33625 ( .A1(n23736), .A2(n23735), .ZN(n23887) );
OR2_X4 U33626 ( .A1(n23737), .A2(n23887), .ZN(n23739) );
NAND2_X4 U33627 ( .A1(n23887), .A2(n23737), .ZN(n23738) );
NAND2_X4 U33628 ( .A1(n23739), .A2(n23738), .ZN(n23879) );
NAND2_X4 U33629 ( .A1(n23740), .A2(n20611), .ZN(n23742) );
OR2_X4 U33630 ( .A1(n20611), .A2(n23740), .ZN(n23741) );
NAND2_X4 U33631 ( .A1(n23742), .A2(n23741), .ZN(n23872) );
NAND2_X4 U33632 ( .A1(n23743), .A2(n20573), .ZN(n23745) );
OR2_X4 U33633 ( .A1(n20573), .A2(n23743), .ZN(n23744) );
NAND2_X4 U33634 ( .A1(n23745), .A2(n23744), .ZN(n23863) );
NAND2_X4 U33635 ( .A1(n23746), .A2(n20535), .ZN(n23748) );
OR2_X4 U33636 ( .A1(n20535), .A2(n23746), .ZN(n23747) );
NAND2_X4 U33637 ( .A1(n23748), .A2(n23747), .ZN(n23856) );
NAND2_X4 U33638 ( .A1(n23749), .A2(n20497), .ZN(n23751) );
OR2_X4 U33639 ( .A1(n20497), .A2(n23749), .ZN(n23750) );
NAND2_X4 U33640 ( .A1(n23751), .A2(n23750), .ZN(n23847) );
NAND2_X4 U33641 ( .A1(n23752), .A2(n20459), .ZN(n23754) );
OR2_X4 U33642 ( .A1(n20459), .A2(n23752), .ZN(n23753) );
NAND2_X4 U33643 ( .A1(n23754), .A2(n23753), .ZN(n23840) );
NAND2_X4 U33644 ( .A1(n23755), .A2(n20421), .ZN(n23757) );
OR2_X4 U33645 ( .A1(n20421), .A2(n23755), .ZN(n23756) );
NAND2_X4 U33646 ( .A1(n23757), .A2(n23756), .ZN(n23831) );
NAND2_X4 U33647 ( .A1(n23758), .A2(n20384), .ZN(n23760) );
OR2_X4 U33648 ( .A1(n20384), .A2(n23758), .ZN(n23759) );
NAND2_X4 U33649 ( .A1(n23760), .A2(n23759), .ZN(n23824) );
NAND2_X4 U33650 ( .A1(n23761), .A2(n20347), .ZN(n23763) );
OR2_X4 U33651 ( .A1(n20347), .A2(n23761), .ZN(n23762) );
NAND2_X4 U33652 ( .A1(n23763), .A2(n23762), .ZN(n23815) );
NAND2_X4 U33653 ( .A1(n23764), .A2(n20310), .ZN(n23766) );
OR2_X4 U33654 ( .A1(n20310), .A2(n23764), .ZN(n23765) );
NAND2_X4 U33655 ( .A1(n23766), .A2(n23765), .ZN(n23808) );
NAND2_X4 U33656 ( .A1(n23767), .A2(n20273), .ZN(n23769) );
OR2_X4 U33657 ( .A1(n20273), .A2(n23767), .ZN(n23768) );
NAND2_X4 U33658 ( .A1(n23769), .A2(n23768), .ZN(n23799) );
NAND2_X4 U33659 ( .A1(n23770), .A2(n20237), .ZN(n23772) );
OR2_X4 U33660 ( .A1(n20237), .A2(n23770), .ZN(n23771) );
NAND2_X4 U33661 ( .A1(n23772), .A2(n23771), .ZN(n23792) );
NAND2_X4 U33662 ( .A1(n23773), .A2(n20201), .ZN(n23775) );
OR2_X4 U33663 ( .A1(n20201), .A2(n23773), .ZN(n23774) );
NAND2_X4 U33664 ( .A1(n23775), .A2(n23774), .ZN(n23939) );
NAND2_X4 U33665 ( .A1(n23776), .A2(n16330), .ZN(n23778) );
OR2_X4 U33666 ( .A1(n16330), .A2(n23776), .ZN(n23777) );
AND2_X4 U33667 ( .A1(n23778), .A2(n23777), .ZN(n23950) );
NAND2_X4 U33668 ( .A1(n20109), .A2(n23779), .ZN(n23784) );
NAND2_X4 U33669 ( .A1(n20167), .A2(n23780), .ZN(n23782) );
NAND2_X4 U33670 ( .A1(n23782), .A2(n23781), .ZN(n23783) );
NAND2_X4 U33671 ( .A1(n23784), .A2(n23783), .ZN(n23949) );
NOR2_X4 U33672 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_0), .ZN(n23948) );
NOR2_X4 U33673 ( .A1(n23949), .A2(n23948), .ZN(n23785) );
OR2_X4 U33674 ( .A1(n23950), .A2(n23785), .ZN(n23787) );
NAND2_X4 U33675 ( .A1(n23785), .A2(n23950), .ZN(n23786) );
NAND2_X4 U33676 ( .A1(n23787), .A2(n23786), .ZN(n25243) );
NAND2_X4 U33677 ( .A1(n25191), .A2(n20083), .ZN(n23790) );
NOR2_X4 U33678 ( .A1(n20762), .A2(n20084), .ZN(n25192) );
NAND2_X4 U33679 ( .A1(n20762), .A2(n20084), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_31_) );
NAND2_X4 U33680 ( .A1(n20081), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_31_), .ZN(n23788) );
NAND2_X4 U33681 ( .A1(n25243), .A2(n23788), .ZN(n23789) );
NAND2_X4 U33682 ( .A1(n23790), .A2(n23789), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N51) );
NAND2_X4 U33683 ( .A1(n20166), .A2(n20201), .ZN(n23796) );
NAND2_X4 U33684 ( .A1(n23792), .A2(n23791), .ZN(n23794) );
NAND2_X4 U33685 ( .A1(n23794), .A2(n23793), .ZN(n23795) );
NAND2_X4 U33686 ( .A1(n23796), .A2(n23795), .ZN(n24100) );
NAND2_X4 U33687 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n24099) );
OR2_X4 U33688 ( .A1(n24100), .A2(n20105), .ZN(n23798) );
NAND2_X4 U33689 ( .A1(n20105), .A2(n24100), .ZN(n23797) );
NAND2_X4 U33690 ( .A1(n23798), .A2(n23797), .ZN(n23936) );
NAND2_X4 U33691 ( .A1(n20202), .A2(n23799), .ZN(n23804) );
NAND2_X4 U33692 ( .A1(n20237), .A2(n23800), .ZN(n23802) );
NAND2_X4 U33693 ( .A1(n23802), .A2(n23801), .ZN(n23803) );
NAND2_X4 U33694 ( .A1(n23804), .A2(n23803), .ZN(n23958) );
NAND2_X4 U33695 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n23956) );
OR2_X4 U33696 ( .A1(n23958), .A2(n20164), .ZN(n23806) );
NAND2_X4 U33697 ( .A1(n20164), .A2(n23958), .ZN(n23805) );
NAND2_X4 U33698 ( .A1(n23806), .A2(n23805), .ZN(n23933) );
NAND2_X4 U33699 ( .A1(n20238), .A2(n20273), .ZN(n23812) );
NAND2_X4 U33700 ( .A1(n23808), .A2(n23807), .ZN(n23810) );
NAND2_X4 U33701 ( .A1(n23810), .A2(n23809), .ZN(n23811) );
NAND2_X4 U33702 ( .A1(n23812), .A2(n23811), .ZN(n23966) );
NAND2_X4 U33703 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n23965) );
OR2_X4 U33704 ( .A1(n23966), .A2(n20200), .ZN(n23814) );
NAND2_X4 U33705 ( .A1(n20200), .A2(n23966), .ZN(n23813) );
NAND2_X4 U33706 ( .A1(n23814), .A2(n23813), .ZN(n23930) );
NAND2_X4 U33707 ( .A1(n20274), .A2(n23815), .ZN(n23820) );
NAND2_X4 U33708 ( .A1(n20310), .A2(n23816), .ZN(n23818) );
NAND2_X4 U33709 ( .A1(n23818), .A2(n23817), .ZN(n23819) );
NAND2_X4 U33710 ( .A1(n23820), .A2(n23819), .ZN(n23974) );
NAND2_X4 U33711 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n23972) );
OR2_X4 U33712 ( .A1(n23974), .A2(n20236), .ZN(n23822) );
NAND2_X4 U33713 ( .A1(n20236), .A2(n23974), .ZN(n23821) );
NAND2_X4 U33714 ( .A1(n23822), .A2(n23821), .ZN(n23927) );
NAND2_X4 U33715 ( .A1(n20311), .A2(n20347), .ZN(n23828) );
NAND2_X4 U33716 ( .A1(n23824), .A2(n23823), .ZN(n23826) );
NAND2_X4 U33717 ( .A1(n23826), .A2(n23825), .ZN(n23827) );
NAND2_X4 U33718 ( .A1(n23828), .A2(n23827), .ZN(n23982) );
NAND2_X4 U33719 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n23981) );
OR2_X4 U33720 ( .A1(n23982), .A2(n20272), .ZN(n23830) );
NAND2_X4 U33721 ( .A1(n20272), .A2(n23982), .ZN(n23829) );
NAND2_X4 U33722 ( .A1(n23830), .A2(n23829), .ZN(n23924) );
NAND2_X4 U33723 ( .A1(n20348), .A2(n23831), .ZN(n23836) );
NAND2_X4 U33724 ( .A1(n20384), .A2(n23832), .ZN(n23834) );
NAND2_X4 U33725 ( .A1(n23834), .A2(n23833), .ZN(n23835) );
NAND2_X4 U33726 ( .A1(n23836), .A2(n23835), .ZN(n23990) );
NAND2_X4 U33727 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n23988) );
OR2_X4 U33728 ( .A1(n23990), .A2(n20309), .ZN(n23838) );
NAND2_X4 U33729 ( .A1(n20309), .A2(n23990), .ZN(n23837) );
NAND2_X4 U33730 ( .A1(n23838), .A2(n23837), .ZN(n23921) );
NAND2_X4 U33731 ( .A1(n20385), .A2(n20421), .ZN(n23844) );
NAND2_X4 U33732 ( .A1(n23840), .A2(n23839), .ZN(n23842) );
NAND2_X4 U33733 ( .A1(n23842), .A2(n23841), .ZN(n23843) );
NAND2_X4 U33734 ( .A1(n23844), .A2(n23843), .ZN(n23998) );
NAND2_X4 U33735 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n23997) );
OR2_X4 U33736 ( .A1(n23998), .A2(n20346), .ZN(n23846) );
NAND2_X4 U33737 ( .A1(n20346), .A2(n23998), .ZN(n23845) );
NAND2_X4 U33738 ( .A1(n23846), .A2(n23845), .ZN(n23918) );
NAND2_X4 U33739 ( .A1(n20422), .A2(n23847), .ZN(n23852) );
NAND2_X4 U33740 ( .A1(n20459), .A2(n23848), .ZN(n23850) );
NAND2_X4 U33741 ( .A1(n23850), .A2(n23849), .ZN(n23851) );
NAND2_X4 U33742 ( .A1(n23852), .A2(n23851), .ZN(n24006) );
NAND2_X4 U33743 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n24004) );
OR2_X4 U33744 ( .A1(n24006), .A2(n20383), .ZN(n23854) );
NAND2_X4 U33745 ( .A1(n20383), .A2(n24006), .ZN(n23853) );
NAND2_X4 U33746 ( .A1(n23854), .A2(n23853), .ZN(n23915) );
NAND2_X4 U33747 ( .A1(n20460), .A2(n20497), .ZN(n23860) );
NAND2_X4 U33748 ( .A1(n23856), .A2(n23855), .ZN(n23858) );
NAND2_X4 U33749 ( .A1(n23858), .A2(n23857), .ZN(n23859) );
NAND2_X4 U33750 ( .A1(n23860), .A2(n23859), .ZN(n24014) );
NAND2_X4 U33751 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n24013) );
OR2_X4 U33752 ( .A1(n24014), .A2(n20420), .ZN(n23862) );
NAND2_X4 U33753 ( .A1(n20420), .A2(n24014), .ZN(n23861) );
NAND2_X4 U33754 ( .A1(n23862), .A2(n23861), .ZN(n23912) );
NAND2_X4 U33755 ( .A1(n20498), .A2(n23863), .ZN(n23868) );
NAND2_X4 U33756 ( .A1(n20535), .A2(n23864), .ZN(n23866) );
NAND2_X4 U33757 ( .A1(n23866), .A2(n23865), .ZN(n23867) );
NAND2_X4 U33758 ( .A1(n23868), .A2(n23867), .ZN(n24022) );
NAND2_X4 U33759 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n24020) );
OR2_X4 U33760 ( .A1(n24022), .A2(n20458), .ZN(n23870) );
NAND2_X4 U33761 ( .A1(n20458), .A2(n24022), .ZN(n23869) );
NAND2_X4 U33762 ( .A1(n23870), .A2(n23869), .ZN(n23909) );
NAND2_X4 U33763 ( .A1(n20536), .A2(n20573), .ZN(n23876) );
NAND2_X4 U33764 ( .A1(n23872), .A2(n23871), .ZN(n23874) );
NAND2_X4 U33765 ( .A1(n23874), .A2(n23873), .ZN(n23875) );
NAND2_X4 U33766 ( .A1(n23876), .A2(n23875), .ZN(n24030) );
NAND2_X4 U33767 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n24029) );
OR2_X4 U33768 ( .A1(n24030), .A2(n20496), .ZN(n23878) );
NAND2_X4 U33769 ( .A1(n20496), .A2(n24030), .ZN(n23877) );
NAND2_X4 U33770 ( .A1(n23878), .A2(n23877), .ZN(n23906) );
NAND2_X4 U33771 ( .A1(n20574), .A2(n23879), .ZN(n23884) );
NAND2_X4 U33772 ( .A1(n20611), .A2(n23880), .ZN(n23882) );
NAND2_X4 U33773 ( .A1(n23882), .A2(n23881), .ZN(n23883) );
NAND2_X4 U33774 ( .A1(n23884), .A2(n23883), .ZN(n24038) );
NAND2_X4 U33775 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n24036) );
OR2_X4 U33776 ( .A1(n24038), .A2(n20534), .ZN(n23886) );
NAND2_X4 U33777 ( .A1(n20534), .A2(n24038), .ZN(n23885) );
NAND2_X4 U33778 ( .A1(n23886), .A2(n23885), .ZN(n23903) );
NAND2_X4 U33779 ( .A1(n23888), .A2(n23887), .ZN(n23890) );
NAND2_X4 U33780 ( .A1(n23890), .A2(n23889), .ZN(n24046) );
NAND2_X4 U33781 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n24045) );
OR2_X4 U33782 ( .A1(n24046), .A2(n20572), .ZN(n23892) );
NAND2_X4 U33783 ( .A1(n20572), .A2(n24046), .ZN(n23891) );
NAND2_X4 U33784 ( .A1(n23892), .A2(n23891), .ZN(n23900) );
NAND2_X4 U33785 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n24054) );
NAND2_X4 U33786 ( .A1(n16200), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_sign_b), .ZN(n23894) );
NOR2_X4 U33787 ( .A1(n23894), .A2(n23893), .ZN(n24056) );
OR2_X4 U33788 ( .A1(n24054), .A2(n24056), .ZN(n23896) );
NAND2_X4 U33789 ( .A1(n24056), .A2(n24054), .ZN(n23895) );
AND2_X4 U33790 ( .A1(n23896), .A2(n23895), .ZN(n23897) );
NOR2_X4 U33791 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_1), .ZN(n24055) );
OR2_X4 U33792 ( .A1(n23897), .A2(n24055), .ZN(n23899) );
NAND2_X4 U33793 ( .A1(n23897), .A2(n24055), .ZN(n23898) );
NAND2_X4 U33794 ( .A1(n23899), .A2(n23898), .ZN(n24044) );
NAND2_X4 U33795 ( .A1(n23900), .A2(n20609), .ZN(n23902) );
OR2_X4 U33796 ( .A1(n20609), .A2(n23900), .ZN(n23901) );
NAND2_X4 U33797 ( .A1(n23902), .A2(n23901), .ZN(n24037) );
NAND2_X4 U33798 ( .A1(n23903), .A2(n20571), .ZN(n23905) );
OR2_X4 U33799 ( .A1(n20571), .A2(n23903), .ZN(n23904) );
NAND2_X4 U33800 ( .A1(n23905), .A2(n23904), .ZN(n24028) );
NAND2_X4 U33801 ( .A1(n23906), .A2(n20533), .ZN(n23908) );
OR2_X4 U33802 ( .A1(n20533), .A2(n23906), .ZN(n23907) );
NAND2_X4 U33803 ( .A1(n23908), .A2(n23907), .ZN(n24021) );
NAND2_X4 U33804 ( .A1(n23909), .A2(n20495), .ZN(n23911) );
OR2_X4 U33805 ( .A1(n20495), .A2(n23909), .ZN(n23910) );
NAND2_X4 U33806 ( .A1(n23911), .A2(n23910), .ZN(n24012) );
NAND2_X4 U33807 ( .A1(n23912), .A2(n20457), .ZN(n23914) );
OR2_X4 U33808 ( .A1(n20457), .A2(n23912), .ZN(n23913) );
NAND2_X4 U33809 ( .A1(n23914), .A2(n23913), .ZN(n24005) );
NAND2_X4 U33810 ( .A1(n23915), .A2(n20419), .ZN(n23917) );
OR2_X4 U33811 ( .A1(n20419), .A2(n23915), .ZN(n23916) );
NAND2_X4 U33812 ( .A1(n23917), .A2(n23916), .ZN(n23996) );
NAND2_X4 U33813 ( .A1(n23918), .A2(n20382), .ZN(n23920) );
OR2_X4 U33814 ( .A1(n20382), .A2(n23918), .ZN(n23919) );
NAND2_X4 U33815 ( .A1(n23920), .A2(n23919), .ZN(n23989) );
NAND2_X4 U33816 ( .A1(n23921), .A2(n20345), .ZN(n23923) );
OR2_X4 U33817 ( .A1(n20345), .A2(n23921), .ZN(n23922) );
NAND2_X4 U33818 ( .A1(n23923), .A2(n23922), .ZN(n23980) );
NAND2_X4 U33819 ( .A1(n23924), .A2(n20308), .ZN(n23926) );
OR2_X4 U33820 ( .A1(n20308), .A2(n23924), .ZN(n23925) );
NAND2_X4 U33821 ( .A1(n23926), .A2(n23925), .ZN(n23973) );
NAND2_X4 U33822 ( .A1(n23927), .A2(n20271), .ZN(n23929) );
OR2_X4 U33823 ( .A1(n20271), .A2(n23927), .ZN(n23928) );
NAND2_X4 U33824 ( .A1(n23929), .A2(n23928), .ZN(n23964) );
NAND2_X4 U33825 ( .A1(n23930), .A2(n20235), .ZN(n23932) );
OR2_X4 U33826 ( .A1(n20235), .A2(n23930), .ZN(n23931) );
NAND2_X4 U33827 ( .A1(n23932), .A2(n23931), .ZN(n23957) );
NAND2_X4 U33828 ( .A1(n23933), .A2(n20199), .ZN(n23935) );
OR2_X4 U33829 ( .A1(n20199), .A2(n23933), .ZN(n23934) );
NAND2_X4 U33830 ( .A1(n23935), .A2(n23934), .ZN(n24098) );
NAND2_X4 U33831 ( .A1(n23936), .A2(n20163), .ZN(n23938) );
OR2_X4 U33832 ( .A1(n20163), .A2(n23936), .ZN(n23937) );
AND2_X4 U33833 ( .A1(n23938), .A2(n23937), .ZN(n24109) );
NAND2_X4 U33834 ( .A1(n20106), .A2(n23939), .ZN(n23944) );
NAND2_X4 U33835 ( .A1(n20165), .A2(n23940), .ZN(n23942) );
NAND2_X4 U33836 ( .A1(n23942), .A2(n23941), .ZN(n23943) );
NAND2_X4 U33837 ( .A1(n23944), .A2(n23943), .ZN(n24108) );
NOR2_X4 U33838 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .ZN(n24107) );
NOR2_X4 U33839 ( .A1(n24108), .A2(n24107), .ZN(n23945) );
OR2_X4 U33840 ( .A1(n24109), .A2(n23945), .ZN(n23947) );
NAND2_X4 U33841 ( .A1(n23945), .A2(n24109), .ZN(n23946) );
NAND2_X4 U33842 ( .A1(n23947), .A2(n23946), .ZN(n23954) );
NAND2_X4 U33843 ( .A1(n23948), .A2(n23950), .ZN(n23952) );
NAND2_X4 U33844 ( .A1(n23950), .A2(n23949), .ZN(n23951) );
NAND2_X4 U33845 ( .A1(n23952), .A2(n23951), .ZN(n23953) );
NOR2_X4 U33846 ( .A1(n23954), .A2(n23953), .ZN(n23955) );
NOR2_X4 U33847 ( .A1(n20082), .A2(n20079), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_16_) );
NOR2_X4 U33848 ( .A1(n23955), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_16_), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_15_) );
NAND2_X4 U33849 ( .A1(n20164), .A2(n20199), .ZN(n23961) );
NAND2_X4 U33850 ( .A1(n23957), .A2(n23956), .ZN(n23959) );
NAND2_X4 U33851 ( .A1(n23959), .A2(n23958), .ZN(n23960) );
NAND2_X4 U33852 ( .A1(n23961), .A2(n23960), .ZN(n24248) );
NAND2_X4 U33853 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n24247) );
OR2_X4 U33854 ( .A1(n24248), .A2(n20104), .ZN(n23963) );
NAND2_X4 U33855 ( .A1(n20104), .A2(n24248), .ZN(n23962) );
NAND2_X4 U33856 ( .A1(n23963), .A2(n23962), .ZN(n24095) );
NAND2_X4 U33857 ( .A1(n20200), .A2(n23964), .ZN(n23969) );
NAND2_X4 U33858 ( .A1(n20235), .A2(n23965), .ZN(n23967) );
NAND2_X4 U33859 ( .A1(n23967), .A2(n23966), .ZN(n23968) );
NAND2_X4 U33860 ( .A1(n23969), .A2(n23968), .ZN(n24117) );
NAND2_X4 U33861 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n24115) );
OR2_X4 U33862 ( .A1(n24117), .A2(n20162), .ZN(n23971) );
NAND2_X4 U33863 ( .A1(n20162), .A2(n24117), .ZN(n23970) );
NAND2_X4 U33864 ( .A1(n23971), .A2(n23970), .ZN(n24092) );
NAND2_X4 U33865 ( .A1(n20236), .A2(n20271), .ZN(n23977) );
NAND2_X4 U33866 ( .A1(n23973), .A2(n23972), .ZN(n23975) );
NAND2_X4 U33867 ( .A1(n23975), .A2(n23974), .ZN(n23976) );
NAND2_X4 U33868 ( .A1(n23977), .A2(n23976), .ZN(n24125) );
NAND2_X4 U33869 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n24124) );
OR2_X4 U33870 ( .A1(n24125), .A2(n20198), .ZN(n23979) );
NAND2_X4 U33871 ( .A1(n20198), .A2(n24125), .ZN(n23978) );
NAND2_X4 U33872 ( .A1(n23979), .A2(n23978), .ZN(n24089) );
NAND2_X4 U33873 ( .A1(n20272), .A2(n23980), .ZN(n23985) );
NAND2_X4 U33874 ( .A1(n20308), .A2(n23981), .ZN(n23983) );
NAND2_X4 U33875 ( .A1(n23983), .A2(n23982), .ZN(n23984) );
NAND2_X4 U33876 ( .A1(n23985), .A2(n23984), .ZN(n24133) );
NAND2_X4 U33877 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n24131) );
OR2_X4 U33878 ( .A1(n24133), .A2(n20234), .ZN(n23987) );
NAND2_X4 U33879 ( .A1(n20234), .A2(n24133), .ZN(n23986) );
NAND2_X4 U33880 ( .A1(n23987), .A2(n23986), .ZN(n24086) );
NAND2_X4 U33881 ( .A1(n20309), .A2(n20345), .ZN(n23993) );
NAND2_X4 U33882 ( .A1(n23989), .A2(n23988), .ZN(n23991) );
NAND2_X4 U33883 ( .A1(n23991), .A2(n23990), .ZN(n23992) );
NAND2_X4 U33884 ( .A1(n23993), .A2(n23992), .ZN(n24141) );
NAND2_X4 U33885 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n24140) );
OR2_X4 U33886 ( .A1(n24141), .A2(n20270), .ZN(n23995) );
NAND2_X4 U33887 ( .A1(n20270), .A2(n24141), .ZN(n23994) );
NAND2_X4 U33888 ( .A1(n23995), .A2(n23994), .ZN(n24083) );
NAND2_X4 U33889 ( .A1(n20346), .A2(n23996), .ZN(n24001) );
NAND2_X4 U33890 ( .A1(n20382), .A2(n23997), .ZN(n23999) );
NAND2_X4 U33891 ( .A1(n23999), .A2(n23998), .ZN(n24000) );
NAND2_X4 U33892 ( .A1(n24001), .A2(n24000), .ZN(n24149) );
NAND2_X4 U33893 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n24147) );
OR2_X4 U33894 ( .A1(n24149), .A2(n20307), .ZN(n24003) );
NAND2_X4 U33895 ( .A1(n20307), .A2(n24149), .ZN(n24002) );
NAND2_X4 U33896 ( .A1(n24003), .A2(n24002), .ZN(n24080) );
NAND2_X4 U33897 ( .A1(n20383), .A2(n20419), .ZN(n24009) );
NAND2_X4 U33898 ( .A1(n24005), .A2(n24004), .ZN(n24007) );
NAND2_X4 U33899 ( .A1(n24007), .A2(n24006), .ZN(n24008) );
NAND2_X4 U33900 ( .A1(n24009), .A2(n24008), .ZN(n24157) );
NAND2_X4 U33901 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n24156) );
OR2_X4 U33902 ( .A1(n24157), .A2(n20344), .ZN(n24011) );
NAND2_X4 U33903 ( .A1(n20344), .A2(n24157), .ZN(n24010) );
NAND2_X4 U33904 ( .A1(n24011), .A2(n24010), .ZN(n24077) );
NAND2_X4 U33905 ( .A1(n20420), .A2(n24012), .ZN(n24017) );
NAND2_X4 U33906 ( .A1(n20457), .A2(n24013), .ZN(n24015) );
NAND2_X4 U33907 ( .A1(n24015), .A2(n24014), .ZN(n24016) );
NAND2_X4 U33908 ( .A1(n24017), .A2(n24016), .ZN(n24165) );
NAND2_X4 U33909 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n24163) );
OR2_X4 U33910 ( .A1(n24165), .A2(n20381), .ZN(n24019) );
NAND2_X4 U33911 ( .A1(n20381), .A2(n24165), .ZN(n24018) );
NAND2_X4 U33912 ( .A1(n24019), .A2(n24018), .ZN(n24074) );
NAND2_X4 U33913 ( .A1(n20458), .A2(n20495), .ZN(n24025) );
NAND2_X4 U33914 ( .A1(n24021), .A2(n24020), .ZN(n24023) );
NAND2_X4 U33915 ( .A1(n24023), .A2(n24022), .ZN(n24024) );
NAND2_X4 U33916 ( .A1(n24025), .A2(n24024), .ZN(n24173) );
NAND2_X4 U33917 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n24172) );
OR2_X4 U33918 ( .A1(n24173), .A2(n20418), .ZN(n24027) );
NAND2_X4 U33919 ( .A1(n20418), .A2(n24173), .ZN(n24026) );
NAND2_X4 U33920 ( .A1(n24027), .A2(n24026), .ZN(n24071) );
NAND2_X4 U33921 ( .A1(n20496), .A2(n24028), .ZN(n24033) );
NAND2_X4 U33922 ( .A1(n20533), .A2(n24029), .ZN(n24031) );
NAND2_X4 U33923 ( .A1(n24031), .A2(n24030), .ZN(n24032) );
NAND2_X4 U33924 ( .A1(n24033), .A2(n24032), .ZN(n24181) );
NAND2_X4 U33925 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n24179) );
OR2_X4 U33926 ( .A1(n24181), .A2(n20456), .ZN(n24035) );
NAND2_X4 U33927 ( .A1(n20456), .A2(n24181), .ZN(n24034) );
NAND2_X4 U33928 ( .A1(n24035), .A2(n24034), .ZN(n24068) );
NAND2_X4 U33929 ( .A1(n20534), .A2(n20571), .ZN(n24041) );
NAND2_X4 U33930 ( .A1(n24037), .A2(n24036), .ZN(n24039) );
NAND2_X4 U33931 ( .A1(n24039), .A2(n24038), .ZN(n24040) );
NAND2_X4 U33932 ( .A1(n24041), .A2(n24040), .ZN(n24189) );
NAND2_X4 U33933 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n24188) );
OR2_X4 U33934 ( .A1(n24189), .A2(n20494), .ZN(n24043) );
NAND2_X4 U33935 ( .A1(n20494), .A2(n24189), .ZN(n24042) );
NAND2_X4 U33936 ( .A1(n24043), .A2(n24042), .ZN(n24065) );
NAND2_X4 U33937 ( .A1(n20572), .A2(n24044), .ZN(n24049) );
NAND2_X4 U33938 ( .A1(n20609), .A2(n24045), .ZN(n24047) );
NAND2_X4 U33939 ( .A1(n24047), .A2(n24046), .ZN(n24048) );
NAND2_X4 U33940 ( .A1(n24049), .A2(n24048), .ZN(n24197) );
NAND2_X4 U33941 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n24195) );
OR2_X4 U33942 ( .A1(n24197), .A2(n20532), .ZN(n24051) );
NAND2_X4 U33943 ( .A1(n20532), .A2(n24197), .ZN(n24050) );
NAND2_X4 U33944 ( .A1(n24051), .A2(n24050), .ZN(n24062) );
NOR2_X4 U33945 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_2), .ZN(n24206) );
NAND2_X4 U33946 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n24205) );
NAND2_X4 U33947 ( .A1(n24206), .A2(n24205), .ZN(n24053) );
OR2_X4 U33948 ( .A1(n24205), .A2(n24206), .ZN(n24052) );
NAND2_X4 U33949 ( .A1(n24053), .A2(n24052), .ZN(n24059) );
NAND2_X4 U33950 ( .A1(n24055), .A2(n20610), .ZN(n24058) );
NAND2_X4 U33951 ( .A1(n20610), .A2(n24056), .ZN(n24057) );
NAND2_X4 U33952 ( .A1(n24058), .A2(n24057), .ZN(n24207) );
NAND2_X4 U33953 ( .A1(n24059), .A2(n24207), .ZN(n24061) );
OR2_X4 U33954 ( .A1(n24207), .A2(n24059), .ZN(n24060) );
NAND2_X4 U33955 ( .A1(n24061), .A2(n24060), .ZN(n24196) );
NAND2_X4 U33956 ( .A1(n24062), .A2(n20569), .ZN(n24064) );
OR2_X4 U33957 ( .A1(n20569), .A2(n24062), .ZN(n24063) );
NAND2_X4 U33958 ( .A1(n24064), .A2(n24063), .ZN(n24187) );
NAND2_X4 U33959 ( .A1(n24065), .A2(n20531), .ZN(n24067) );
OR2_X4 U33960 ( .A1(n20531), .A2(n24065), .ZN(n24066) );
NAND2_X4 U33961 ( .A1(n24067), .A2(n24066), .ZN(n24180) );
NAND2_X4 U33962 ( .A1(n24068), .A2(n20493), .ZN(n24070) );
OR2_X4 U33963 ( .A1(n20493), .A2(n24068), .ZN(n24069) );
NAND2_X4 U33964 ( .A1(n24070), .A2(n24069), .ZN(n24171) );
NAND2_X4 U33965 ( .A1(n24071), .A2(n20455), .ZN(n24073) );
OR2_X4 U33966 ( .A1(n20455), .A2(n24071), .ZN(n24072) );
NAND2_X4 U33967 ( .A1(n24073), .A2(n24072), .ZN(n24164) );
NAND2_X4 U33968 ( .A1(n24074), .A2(n20417), .ZN(n24076) );
OR2_X4 U33969 ( .A1(n20417), .A2(n24074), .ZN(n24075) );
NAND2_X4 U33970 ( .A1(n24076), .A2(n24075), .ZN(n24155) );
NAND2_X4 U33971 ( .A1(n24077), .A2(n20380), .ZN(n24079) );
OR2_X4 U33972 ( .A1(n20380), .A2(n24077), .ZN(n24078) );
NAND2_X4 U33973 ( .A1(n24079), .A2(n24078), .ZN(n24148) );
NAND2_X4 U33974 ( .A1(n24080), .A2(n20343), .ZN(n24082) );
OR2_X4 U33975 ( .A1(n20343), .A2(n24080), .ZN(n24081) );
NAND2_X4 U33976 ( .A1(n24082), .A2(n24081), .ZN(n24139) );
NAND2_X4 U33977 ( .A1(n24083), .A2(n20306), .ZN(n24085) );
OR2_X4 U33978 ( .A1(n20306), .A2(n24083), .ZN(n24084) );
NAND2_X4 U33979 ( .A1(n24085), .A2(n24084), .ZN(n24132) );
NAND2_X4 U33980 ( .A1(n24086), .A2(n20269), .ZN(n24088) );
OR2_X4 U33981 ( .A1(n20269), .A2(n24086), .ZN(n24087) );
NAND2_X4 U33982 ( .A1(n24088), .A2(n24087), .ZN(n24123) );
NAND2_X4 U33983 ( .A1(n24089), .A2(n20233), .ZN(n24091) );
OR2_X4 U33984 ( .A1(n20233), .A2(n24089), .ZN(n24090) );
NAND2_X4 U33985 ( .A1(n24091), .A2(n24090), .ZN(n24116) );
NAND2_X4 U33986 ( .A1(n24092), .A2(n20197), .ZN(n24094) );
OR2_X4 U33987 ( .A1(n20197), .A2(n24092), .ZN(n24093) );
NAND2_X4 U33988 ( .A1(n24094), .A2(n24093), .ZN(n24246) );
NAND2_X4 U33989 ( .A1(n24095), .A2(n20161), .ZN(n24097) );
OR2_X4 U33990 ( .A1(n20161), .A2(n24095), .ZN(n24096) );
AND2_X4 U33991 ( .A1(n24097), .A2(n24096), .ZN(n24257) );
NAND2_X4 U33992 ( .A1(n20105), .A2(n24098), .ZN(n24103) );
NAND2_X4 U33993 ( .A1(n20163), .A2(n24099), .ZN(n24101) );
NAND2_X4 U33994 ( .A1(n24101), .A2(n24100), .ZN(n24102) );
NAND2_X4 U33995 ( .A1(n24103), .A2(n24102), .ZN(n24256) );
NOR2_X4 U33996 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_2), .ZN(n24255) );
NOR2_X4 U33997 ( .A1(n24256), .A2(n24255), .ZN(n24104) );
OR2_X4 U33998 ( .A1(n24257), .A2(n24104), .ZN(n24106) );
NAND2_X4 U33999 ( .A1(n24104), .A2(n24257), .ZN(n24105) );
NAND2_X4 U34000 ( .A1(n24106), .A2(n24105), .ZN(n24113) );
NAND2_X4 U34001 ( .A1(n24107), .A2(n24109), .ZN(n24111) );
NAND2_X4 U34002 ( .A1(n24109), .A2(n24108), .ZN(n24110) );
NAND2_X4 U34003 ( .A1(n24111), .A2(n24110), .ZN(n24112) );
NOR2_X4 U34004 ( .A1(n24113), .A2(n24112), .ZN(n24114) );
NOR2_X4 U34005 ( .A1(n20077), .A2(n20076), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_17_) );
NOR2_X4 U34006 ( .A1(n24114), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_17_), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_16_) );
NAND2_X4 U34007 ( .A1(n20162), .A2(n20197), .ZN(n24120) );
NAND2_X4 U34008 ( .A1(n24116), .A2(n24115), .ZN(n24118) );
NAND2_X4 U34009 ( .A1(n24118), .A2(n24117), .ZN(n24119) );
NAND2_X4 U34010 ( .A1(n24120), .A2(n24119), .ZN(n24384) );
NAND2_X4 U34011 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n24382) );
OR2_X4 U34012 ( .A1(n24384), .A2(n20103), .ZN(n24122) );
NAND2_X4 U34013 ( .A1(n20103), .A2(n24384), .ZN(n24121) );
NAND2_X4 U34014 ( .A1(n24122), .A2(n24121), .ZN(n24243) );
NAND2_X4 U34015 ( .A1(n20198), .A2(n24123), .ZN(n24128) );
NAND2_X4 U34016 ( .A1(n20233), .A2(n24124), .ZN(n24126) );
NAND2_X4 U34017 ( .A1(n24126), .A2(n24125), .ZN(n24127) );
NAND2_X4 U34018 ( .A1(n24128), .A2(n24127), .ZN(n24264) );
NAND2_X4 U34019 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n24263) );
OR2_X4 U34020 ( .A1(n24264), .A2(n20160), .ZN(n24130) );
NAND2_X4 U34021 ( .A1(n20160), .A2(n24264), .ZN(n24129) );
NAND2_X4 U34022 ( .A1(n24130), .A2(n24129), .ZN(n24240) );
NAND2_X4 U34023 ( .A1(n20234), .A2(n20269), .ZN(n24136) );
NAND2_X4 U34024 ( .A1(n24132), .A2(n24131), .ZN(n24134) );
NAND2_X4 U34025 ( .A1(n24134), .A2(n24133), .ZN(n24135) );
NAND2_X4 U34026 ( .A1(n24136), .A2(n24135), .ZN(n24272) );
NAND2_X4 U34027 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n24270) );
OR2_X4 U34028 ( .A1(n24272), .A2(n20196), .ZN(n24138) );
NAND2_X4 U34029 ( .A1(n20196), .A2(n24272), .ZN(n24137) );
NAND2_X4 U34030 ( .A1(n24138), .A2(n24137), .ZN(n24237) );
NAND2_X4 U34031 ( .A1(n20270), .A2(n24139), .ZN(n24144) );
NAND2_X4 U34032 ( .A1(n20306), .A2(n24140), .ZN(n24142) );
NAND2_X4 U34033 ( .A1(n24142), .A2(n24141), .ZN(n24143) );
NAND2_X4 U34034 ( .A1(n24144), .A2(n24143), .ZN(n24280) );
NAND2_X4 U34035 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n24279) );
OR2_X4 U34036 ( .A1(n24280), .A2(n20232), .ZN(n24146) );
NAND2_X4 U34037 ( .A1(n20232), .A2(n24280), .ZN(n24145) );
NAND2_X4 U34038 ( .A1(n24146), .A2(n24145), .ZN(n24234) );
NAND2_X4 U34039 ( .A1(n20307), .A2(n20343), .ZN(n24152) );
NAND2_X4 U34040 ( .A1(n24148), .A2(n24147), .ZN(n24150) );
NAND2_X4 U34041 ( .A1(n24150), .A2(n24149), .ZN(n24151) );
NAND2_X4 U34042 ( .A1(n24152), .A2(n24151), .ZN(n24288) );
NAND2_X4 U34043 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n24286) );
OR2_X4 U34044 ( .A1(n24288), .A2(n20268), .ZN(n24154) );
NAND2_X4 U34045 ( .A1(n20268), .A2(n24288), .ZN(n24153) );
NAND2_X4 U34046 ( .A1(n24154), .A2(n24153), .ZN(n24231) );
NAND2_X4 U34047 ( .A1(n20344), .A2(n24155), .ZN(n24160) );
NAND2_X4 U34048 ( .A1(n20380), .A2(n24156), .ZN(n24158) );
NAND2_X4 U34049 ( .A1(n24158), .A2(n24157), .ZN(n24159) );
NAND2_X4 U34050 ( .A1(n24160), .A2(n24159), .ZN(n24296) );
NAND2_X4 U34051 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n24295) );
OR2_X4 U34052 ( .A1(n24296), .A2(n20305), .ZN(n24162) );
NAND2_X4 U34053 ( .A1(n20305), .A2(n24296), .ZN(n24161) );
NAND2_X4 U34054 ( .A1(n24162), .A2(n24161), .ZN(n24228) );
NAND2_X4 U34055 ( .A1(n20381), .A2(n20417), .ZN(n24168) );
NAND2_X4 U34056 ( .A1(n24164), .A2(n24163), .ZN(n24166) );
NAND2_X4 U34057 ( .A1(n24166), .A2(n24165), .ZN(n24167) );
NAND2_X4 U34058 ( .A1(n24168), .A2(n24167), .ZN(n24304) );
NAND2_X4 U34059 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n24302) );
OR2_X4 U34060 ( .A1(n24304), .A2(n20342), .ZN(n24170) );
NAND2_X4 U34061 ( .A1(n20342), .A2(n24304), .ZN(n24169) );
NAND2_X4 U34062 ( .A1(n24170), .A2(n24169), .ZN(n24225) );
NAND2_X4 U34063 ( .A1(n20418), .A2(n24171), .ZN(n24176) );
NAND2_X4 U34064 ( .A1(n20455), .A2(n24172), .ZN(n24174) );
NAND2_X4 U34065 ( .A1(n24174), .A2(n24173), .ZN(n24175) );
NAND2_X4 U34066 ( .A1(n24176), .A2(n24175), .ZN(n24312) );
NAND2_X4 U34067 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n24311) );
OR2_X4 U34068 ( .A1(n24312), .A2(n20379), .ZN(n24178) );
NAND2_X4 U34069 ( .A1(n20379), .A2(n24312), .ZN(n24177) );
NAND2_X4 U34070 ( .A1(n24178), .A2(n24177), .ZN(n24222) );
NAND2_X4 U34071 ( .A1(n20456), .A2(n20493), .ZN(n24184) );
NAND2_X4 U34072 ( .A1(n24180), .A2(n24179), .ZN(n24182) );
NAND2_X4 U34073 ( .A1(n24182), .A2(n24181), .ZN(n24183) );
NAND2_X4 U34074 ( .A1(n24184), .A2(n24183), .ZN(n24320) );
NAND2_X4 U34075 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n24318) );
OR2_X4 U34076 ( .A1(n24320), .A2(n20416), .ZN(n24186) );
NAND2_X4 U34077 ( .A1(n20416), .A2(n24320), .ZN(n24185) );
NAND2_X4 U34078 ( .A1(n24186), .A2(n24185), .ZN(n24219) );
NAND2_X4 U34079 ( .A1(n20494), .A2(n24187), .ZN(n24192) );
NAND2_X4 U34080 ( .A1(n20531), .A2(n24188), .ZN(n24190) );
NAND2_X4 U34081 ( .A1(n24190), .A2(n24189), .ZN(n24191) );
NAND2_X4 U34082 ( .A1(n24192), .A2(n24191), .ZN(n24328) );
NAND2_X4 U34083 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n24327) );
OR2_X4 U34084 ( .A1(n24328), .A2(n20454), .ZN(n24194) );
NAND2_X4 U34085 ( .A1(n20454), .A2(n24328), .ZN(n24193) );
NAND2_X4 U34086 ( .A1(n24194), .A2(n24193), .ZN(n24216) );
NAND2_X4 U34087 ( .A1(n20532), .A2(n20569), .ZN(n24200) );
NAND2_X4 U34088 ( .A1(n24196), .A2(n24195), .ZN(n24198) );
NAND2_X4 U34089 ( .A1(n24198), .A2(n24197), .ZN(n24199) );
NAND2_X4 U34090 ( .A1(n24200), .A2(n24199), .ZN(n24336) );
NAND2_X4 U34091 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n24334) );
OR2_X4 U34092 ( .A1(n24336), .A2(n20492), .ZN(n24202) );
NAND2_X4 U34093 ( .A1(n20492), .A2(n24336), .ZN(n24201) );
NAND2_X4 U34094 ( .A1(n24202), .A2(n24201), .ZN(n24213) );
NOR2_X4 U34095 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_3), .ZN(n24345) );
NAND2_X4 U34096 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n24344) );
NAND2_X4 U34097 ( .A1(n24345), .A2(n24344), .ZN(n24204) );
OR2_X4 U34098 ( .A1(n24344), .A2(n24345), .ZN(n24203) );
NAND2_X4 U34099 ( .A1(n24204), .A2(n24203), .ZN(n24210) );
NAND2_X4 U34100 ( .A1(n24206), .A2(n20570), .ZN(n24209) );
NAND2_X4 U34101 ( .A1(n20570), .A2(n24207), .ZN(n24208) );
NAND2_X4 U34102 ( .A1(n24209), .A2(n24208), .ZN(n24346) );
NAND2_X4 U34103 ( .A1(n24210), .A2(n24346), .ZN(n24212) );
OR2_X4 U34104 ( .A1(n24346), .A2(n24210), .ZN(n24211) );
NAND2_X4 U34105 ( .A1(n24212), .A2(n24211), .ZN(n24335) );
NAND2_X4 U34106 ( .A1(n24213), .A2(n20529), .ZN(n24215) );
OR2_X4 U34107 ( .A1(n20529), .A2(n24213), .ZN(n24214) );
NAND2_X4 U34108 ( .A1(n24215), .A2(n24214), .ZN(n24326) );
NAND2_X4 U34109 ( .A1(n24216), .A2(n20491), .ZN(n24218) );
OR2_X4 U34110 ( .A1(n20491), .A2(n24216), .ZN(n24217) );
NAND2_X4 U34111 ( .A1(n24218), .A2(n24217), .ZN(n24319) );
NAND2_X4 U34112 ( .A1(n24219), .A2(n20453), .ZN(n24221) );
OR2_X4 U34113 ( .A1(n20453), .A2(n24219), .ZN(n24220) );
NAND2_X4 U34114 ( .A1(n24221), .A2(n24220), .ZN(n24310) );
NAND2_X4 U34115 ( .A1(n24222), .A2(n20415), .ZN(n24224) );
OR2_X4 U34116 ( .A1(n20415), .A2(n24222), .ZN(n24223) );
NAND2_X4 U34117 ( .A1(n24224), .A2(n24223), .ZN(n24303) );
NAND2_X4 U34118 ( .A1(n24225), .A2(n20378), .ZN(n24227) );
OR2_X4 U34119 ( .A1(n20378), .A2(n24225), .ZN(n24226) );
NAND2_X4 U34120 ( .A1(n24227), .A2(n24226), .ZN(n24294) );
NAND2_X4 U34121 ( .A1(n24228), .A2(n20341), .ZN(n24230) );
OR2_X4 U34122 ( .A1(n20341), .A2(n24228), .ZN(n24229) );
NAND2_X4 U34123 ( .A1(n24230), .A2(n24229), .ZN(n24287) );
NAND2_X4 U34124 ( .A1(n24231), .A2(n20304), .ZN(n24233) );
OR2_X4 U34125 ( .A1(n20304), .A2(n24231), .ZN(n24232) );
NAND2_X4 U34126 ( .A1(n24233), .A2(n24232), .ZN(n24278) );
NAND2_X4 U34127 ( .A1(n24234), .A2(n20267), .ZN(n24236) );
OR2_X4 U34128 ( .A1(n20267), .A2(n24234), .ZN(n24235) );
NAND2_X4 U34129 ( .A1(n24236), .A2(n24235), .ZN(n24271) );
NAND2_X4 U34130 ( .A1(n24237), .A2(n20231), .ZN(n24239) );
OR2_X4 U34131 ( .A1(n20231), .A2(n24237), .ZN(n24238) );
NAND2_X4 U34132 ( .A1(n24239), .A2(n24238), .ZN(n24262) );
NAND2_X4 U34133 ( .A1(n24240), .A2(n20195), .ZN(n24242) );
OR2_X4 U34134 ( .A1(n20195), .A2(n24240), .ZN(n24241) );
NAND2_X4 U34135 ( .A1(n24242), .A2(n24241), .ZN(n24383) );
NAND2_X4 U34136 ( .A1(n24243), .A2(n20159), .ZN(n24245) );
OR2_X4 U34137 ( .A1(n20159), .A2(n24243), .ZN(n24244) );
NAND2_X4 U34138 ( .A1(n24245), .A2(n24244), .ZN(n24393) );
NAND2_X4 U34139 ( .A1(n20104), .A2(n24246), .ZN(n24251) );
NAND2_X4 U34140 ( .A1(n20161), .A2(n24247), .ZN(n24249) );
NAND2_X4 U34141 ( .A1(n24249), .A2(n24248), .ZN(n24250) );
NAND2_X4 U34142 ( .A1(n24251), .A2(n24250), .ZN(n24392) );
NOR2_X4 U34143 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_3), .ZN(n24391) );
NOR2_X4 U34144 ( .A1(n24392), .A2(n24391), .ZN(n24252) );
OR2_X4 U34145 ( .A1(n20102), .A2(n24252), .ZN(n24254) );
NAND2_X4 U34146 ( .A1(n24252), .A2(n20102), .ZN(n24253) );
NAND2_X4 U34147 ( .A1(n24254), .A2(n24253), .ZN(n25246) );
NAND2_X4 U34148 ( .A1(n24255), .A2(n24257), .ZN(n24259) );
NAND2_X4 U34149 ( .A1(n24257), .A2(n24256), .ZN(n24258) );
NAND2_X4 U34150 ( .A1(n24259), .A2(n24258), .ZN(n25245) );
NAND2_X4 U34151 ( .A1(n25246), .A2(n25245), .ZN(n24261) );
OR2_X4 U34152 ( .A1(n25245), .A2(n25246), .ZN(n24260) );
NAND2_X4 U34153 ( .A1(n24261), .A2(n24260), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_17_) );
NAND2_X4 U34154 ( .A1(n20160), .A2(n24262), .ZN(n24267) );
NAND2_X4 U34155 ( .A1(n20195), .A2(n24263), .ZN(n24265) );
NAND2_X4 U34156 ( .A1(n24265), .A2(n24264), .ZN(n24266) );
NAND2_X4 U34157 ( .A1(n24267), .A2(n24266), .ZN(n24510) );
NAND2_X4 U34158 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n24509) );
OR2_X4 U34159 ( .A1(n24510), .A2(n20101), .ZN(n24269) );
NAND2_X4 U34160 ( .A1(n20101), .A2(n24510), .ZN(n24268) );
NAND2_X4 U34161 ( .A1(n24269), .A2(n24268), .ZN(n24379) );
NAND2_X4 U34162 ( .A1(n20196), .A2(n20231), .ZN(n24275) );
NAND2_X4 U34163 ( .A1(n24271), .A2(n24270), .ZN(n24273) );
NAND2_X4 U34164 ( .A1(n24273), .A2(n24272), .ZN(n24274) );
NAND2_X4 U34165 ( .A1(n24275), .A2(n24274), .ZN(n24401) );
NAND2_X4 U34166 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n24399) );
OR2_X4 U34167 ( .A1(n24401), .A2(n20158), .ZN(n24277) );
NAND2_X4 U34168 ( .A1(n20158), .A2(n24401), .ZN(n24276) );
NAND2_X4 U34169 ( .A1(n24277), .A2(n24276), .ZN(n24376) );
NAND2_X4 U34170 ( .A1(n20232), .A2(n24278), .ZN(n24283) );
NAND2_X4 U34171 ( .A1(n20267), .A2(n24279), .ZN(n24281) );
NAND2_X4 U34172 ( .A1(n24281), .A2(n24280), .ZN(n24282) );
NAND2_X4 U34173 ( .A1(n24283), .A2(n24282), .ZN(n24409) );
NAND2_X4 U34174 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n24408) );
OR2_X4 U34175 ( .A1(n24409), .A2(n20194), .ZN(n24285) );
NAND2_X4 U34176 ( .A1(n20194), .A2(n24409), .ZN(n24284) );
NAND2_X4 U34177 ( .A1(n24285), .A2(n24284), .ZN(n24373) );
NAND2_X4 U34178 ( .A1(n20268), .A2(n20304), .ZN(n24291) );
NAND2_X4 U34179 ( .A1(n24287), .A2(n24286), .ZN(n24289) );
NAND2_X4 U34180 ( .A1(n24289), .A2(n24288), .ZN(n24290) );
NAND2_X4 U34181 ( .A1(n24291), .A2(n24290), .ZN(n24417) );
NAND2_X4 U34182 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n24415) );
OR2_X4 U34183 ( .A1(n24417), .A2(n20230), .ZN(n24293) );
NAND2_X4 U34184 ( .A1(n20230), .A2(n24417), .ZN(n24292) );
NAND2_X4 U34185 ( .A1(n24293), .A2(n24292), .ZN(n24370) );
NAND2_X4 U34186 ( .A1(n20305), .A2(n24294), .ZN(n24299) );
NAND2_X4 U34187 ( .A1(n20341), .A2(n24295), .ZN(n24297) );
NAND2_X4 U34188 ( .A1(n24297), .A2(n24296), .ZN(n24298) );
NAND2_X4 U34189 ( .A1(n24299), .A2(n24298), .ZN(n24425) );
NAND2_X4 U34190 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n24424) );
OR2_X4 U34191 ( .A1(n24425), .A2(n20266), .ZN(n24301) );
NAND2_X4 U34192 ( .A1(n20266), .A2(n24425), .ZN(n24300) );
NAND2_X4 U34193 ( .A1(n24301), .A2(n24300), .ZN(n24367) );
NAND2_X4 U34194 ( .A1(n20342), .A2(n20378), .ZN(n24307) );
NAND2_X4 U34195 ( .A1(n24303), .A2(n24302), .ZN(n24305) );
NAND2_X4 U34196 ( .A1(n24305), .A2(n24304), .ZN(n24306) );
NAND2_X4 U34197 ( .A1(n24307), .A2(n24306), .ZN(n24433) );
NAND2_X4 U34198 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n24431) );
OR2_X4 U34199 ( .A1(n24433), .A2(n20303), .ZN(n24309) );
NAND2_X4 U34200 ( .A1(n20303), .A2(n24433), .ZN(n24308) );
NAND2_X4 U34201 ( .A1(n24309), .A2(n24308), .ZN(n24364) );
NAND2_X4 U34202 ( .A1(n20379), .A2(n24310), .ZN(n24315) );
NAND2_X4 U34203 ( .A1(n20415), .A2(n24311), .ZN(n24313) );
NAND2_X4 U34204 ( .A1(n24313), .A2(n24312), .ZN(n24314) );
NAND2_X4 U34205 ( .A1(n24315), .A2(n24314), .ZN(n24441) );
NAND2_X4 U34206 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n24440) );
OR2_X4 U34207 ( .A1(n24441), .A2(n20340), .ZN(n24317) );
NAND2_X4 U34208 ( .A1(n20340), .A2(n24441), .ZN(n24316) );
NAND2_X4 U34209 ( .A1(n24317), .A2(n24316), .ZN(n24361) );
NAND2_X4 U34210 ( .A1(n20416), .A2(n20453), .ZN(n24323) );
NAND2_X4 U34211 ( .A1(n24319), .A2(n24318), .ZN(n24321) );
NAND2_X4 U34212 ( .A1(n24321), .A2(n24320), .ZN(n24322) );
NAND2_X4 U34213 ( .A1(n24323), .A2(n24322), .ZN(n24449) );
NAND2_X4 U34214 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n24447) );
OR2_X4 U34215 ( .A1(n24449), .A2(n20377), .ZN(n24325) );
NAND2_X4 U34216 ( .A1(n20377), .A2(n24449), .ZN(n24324) );
NAND2_X4 U34217 ( .A1(n24325), .A2(n24324), .ZN(n24358) );
NAND2_X4 U34218 ( .A1(n20454), .A2(n24326), .ZN(n24331) );
NAND2_X4 U34219 ( .A1(n20491), .A2(n24327), .ZN(n24329) );
NAND2_X4 U34220 ( .A1(n24329), .A2(n24328), .ZN(n24330) );
NAND2_X4 U34221 ( .A1(n24331), .A2(n24330), .ZN(n24457) );
NAND2_X4 U34222 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n24456) );
OR2_X4 U34223 ( .A1(n24457), .A2(n20414), .ZN(n24333) );
NAND2_X4 U34224 ( .A1(n20414), .A2(n24457), .ZN(n24332) );
NAND2_X4 U34225 ( .A1(n24333), .A2(n24332), .ZN(n24355) );
NAND2_X4 U34226 ( .A1(n20492), .A2(n20529), .ZN(n24339) );
NAND2_X4 U34227 ( .A1(n24335), .A2(n24334), .ZN(n24337) );
NAND2_X4 U34228 ( .A1(n24337), .A2(n24336), .ZN(n24338) );
NAND2_X4 U34229 ( .A1(n24339), .A2(n24338), .ZN(n24465) );
NAND2_X4 U34230 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n24463) );
OR2_X4 U34231 ( .A1(n24465), .A2(n20452), .ZN(n24341) );
NAND2_X4 U34232 ( .A1(n20452), .A2(n24465), .ZN(n24340) );
NAND2_X4 U34233 ( .A1(n24341), .A2(n24340), .ZN(n24352) );
NOR2_X4 U34234 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_4), .ZN(n24474) );
NAND2_X4 U34235 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n24473) );
NAND2_X4 U34236 ( .A1(n24474), .A2(n24473), .ZN(n24343) );
OR2_X4 U34237 ( .A1(n24473), .A2(n24474), .ZN(n24342) );
NAND2_X4 U34238 ( .A1(n24343), .A2(n24342), .ZN(n24349) );
NAND2_X4 U34239 ( .A1(n24345), .A2(n20530), .ZN(n24348) );
NAND2_X4 U34240 ( .A1(n20530), .A2(n24346), .ZN(n24347) );
NAND2_X4 U34241 ( .A1(n24348), .A2(n24347), .ZN(n24475) );
NAND2_X4 U34242 ( .A1(n24349), .A2(n24475), .ZN(n24351) );
OR2_X4 U34243 ( .A1(n24475), .A2(n24349), .ZN(n24350) );
NAND2_X4 U34244 ( .A1(n24351), .A2(n24350), .ZN(n24464) );
NAND2_X4 U34245 ( .A1(n24352), .A2(n20489), .ZN(n24354) );
OR2_X4 U34246 ( .A1(n20489), .A2(n24352), .ZN(n24353) );
NAND2_X4 U34247 ( .A1(n24354), .A2(n24353), .ZN(n24455) );
NAND2_X4 U34248 ( .A1(n24355), .A2(n20451), .ZN(n24357) );
OR2_X4 U34249 ( .A1(n20451), .A2(n24355), .ZN(n24356) );
NAND2_X4 U34250 ( .A1(n24357), .A2(n24356), .ZN(n24448) );
NAND2_X4 U34251 ( .A1(n24358), .A2(n20413), .ZN(n24360) );
OR2_X4 U34252 ( .A1(n20413), .A2(n24358), .ZN(n24359) );
NAND2_X4 U34253 ( .A1(n24360), .A2(n24359), .ZN(n24439) );
NAND2_X4 U34254 ( .A1(n24361), .A2(n20376), .ZN(n24363) );
OR2_X4 U34255 ( .A1(n20376), .A2(n24361), .ZN(n24362) );
NAND2_X4 U34256 ( .A1(n24363), .A2(n24362), .ZN(n24432) );
NAND2_X4 U34257 ( .A1(n24364), .A2(n20339), .ZN(n24366) );
OR2_X4 U34258 ( .A1(n20339), .A2(n24364), .ZN(n24365) );
NAND2_X4 U34259 ( .A1(n24366), .A2(n24365), .ZN(n24423) );
NAND2_X4 U34260 ( .A1(n24367), .A2(n20302), .ZN(n24369) );
OR2_X4 U34261 ( .A1(n20302), .A2(n24367), .ZN(n24368) );
NAND2_X4 U34262 ( .A1(n24369), .A2(n24368), .ZN(n24416) );
NAND2_X4 U34263 ( .A1(n24370), .A2(n20265), .ZN(n24372) );
OR2_X4 U34264 ( .A1(n20265), .A2(n24370), .ZN(n24371) );
NAND2_X4 U34265 ( .A1(n24372), .A2(n24371), .ZN(n24407) );
NAND2_X4 U34266 ( .A1(n24373), .A2(n20229), .ZN(n24375) );
OR2_X4 U34267 ( .A1(n20229), .A2(n24373), .ZN(n24374) );
NAND2_X4 U34268 ( .A1(n24375), .A2(n24374), .ZN(n24400) );
NAND2_X4 U34269 ( .A1(n24376), .A2(n20193), .ZN(n24378) );
OR2_X4 U34270 ( .A1(n20193), .A2(n24376), .ZN(n24377) );
NAND2_X4 U34271 ( .A1(n24378), .A2(n24377), .ZN(n24508) );
NAND2_X4 U34272 ( .A1(n24379), .A2(n20157), .ZN(n24381) );
OR2_X4 U34273 ( .A1(n20157), .A2(n24379), .ZN(n24380) );
AND2_X4 U34274 ( .A1(n24381), .A2(n24380), .ZN(n24519) );
NAND2_X4 U34275 ( .A1(n20103), .A2(n20159), .ZN(n24387) );
NAND2_X4 U34276 ( .A1(n24383), .A2(n24382), .ZN(n24385) );
NAND2_X4 U34277 ( .A1(n24385), .A2(n24384), .ZN(n24386) );
NAND2_X4 U34278 ( .A1(n24387), .A2(n24386), .ZN(n24518) );
NOR2_X4 U34279 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_4), .ZN(n24517) );
NOR2_X4 U34280 ( .A1(n24518), .A2(n24517), .ZN(n24388) );
OR2_X4 U34281 ( .A1(n24519), .A2(n24388), .ZN(n24390) );
NAND2_X4 U34282 ( .A1(n24388), .A2(n24519), .ZN(n24389) );
NAND2_X4 U34283 ( .A1(n24390), .A2(n24389), .ZN(n24397) );
NAND2_X4 U34284 ( .A1(n24391), .A2(n24393), .ZN(n24395) );
NAND2_X4 U34285 ( .A1(n24393), .A2(n24392), .ZN(n24394) );
NAND2_X4 U34286 ( .A1(n24395), .A2(n24394), .ZN(n24396) );
NOR2_X4 U34287 ( .A1(n24397), .A2(n24396), .ZN(n24398) );
NOR2_X4 U34288 ( .A1(n20070), .A2(n20069), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_19_) );
NOR2_X4 U34289 ( .A1(n24398), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_19_), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_18_) );
NAND2_X4 U34290 ( .A1(n20158), .A2(n20193), .ZN(n24404) );
NAND2_X4 U34291 ( .A1(n24400), .A2(n24399), .ZN(n24402) );
NAND2_X4 U34292 ( .A1(n24402), .A2(n24401), .ZN(n24403) );
NAND2_X4 U34293 ( .A1(n24404), .A2(n24403), .ZN(n24630) );
NAND2_X4 U34294 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n24628) );
OR2_X4 U34295 ( .A1(n24630), .A2(n20100), .ZN(n24406) );
NAND2_X4 U34296 ( .A1(n20100), .A2(n24630), .ZN(n24405) );
NAND2_X4 U34297 ( .A1(n24406), .A2(n24405), .ZN(n24505) );
NAND2_X4 U34298 ( .A1(n20194), .A2(n24407), .ZN(n24412) );
NAND2_X4 U34299 ( .A1(n20229), .A2(n24408), .ZN(n24410) );
NAND2_X4 U34300 ( .A1(n24410), .A2(n24409), .ZN(n24411) );
NAND2_X4 U34301 ( .A1(n24412), .A2(n24411), .ZN(n24532) );
NAND2_X4 U34302 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n24531) );
OR2_X4 U34303 ( .A1(n24532), .A2(n20156), .ZN(n24414) );
NAND2_X4 U34304 ( .A1(n20156), .A2(n24532), .ZN(n24413) );
NAND2_X4 U34305 ( .A1(n24414), .A2(n24413), .ZN(n24502) );
NAND2_X4 U34306 ( .A1(n20230), .A2(n20265), .ZN(n24420) );
NAND2_X4 U34307 ( .A1(n24416), .A2(n24415), .ZN(n24418) );
NAND2_X4 U34308 ( .A1(n24418), .A2(n24417), .ZN(n24419) );
NAND2_X4 U34309 ( .A1(n24420), .A2(n24419), .ZN(n24540) );
NAND2_X4 U34310 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n24538) );
OR2_X4 U34311 ( .A1(n24540), .A2(n20192), .ZN(n24422) );
NAND2_X4 U34312 ( .A1(n20192), .A2(n24540), .ZN(n24421) );
NAND2_X4 U34313 ( .A1(n24422), .A2(n24421), .ZN(n24499) );
NAND2_X4 U34314 ( .A1(n20266), .A2(n24423), .ZN(n24428) );
NAND2_X4 U34315 ( .A1(n20302), .A2(n24424), .ZN(n24426) );
NAND2_X4 U34316 ( .A1(n24426), .A2(n24425), .ZN(n24427) );
NAND2_X4 U34317 ( .A1(n24428), .A2(n24427), .ZN(n24548) );
NAND2_X4 U34318 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n24547) );
OR2_X4 U34319 ( .A1(n24548), .A2(n20228), .ZN(n24430) );
NAND2_X4 U34320 ( .A1(n20228), .A2(n24548), .ZN(n24429) );
NAND2_X4 U34321 ( .A1(n24430), .A2(n24429), .ZN(n24496) );
NAND2_X4 U34322 ( .A1(n20303), .A2(n20339), .ZN(n24436) );
NAND2_X4 U34323 ( .A1(n24432), .A2(n24431), .ZN(n24434) );
NAND2_X4 U34324 ( .A1(n24434), .A2(n24433), .ZN(n24435) );
NAND2_X4 U34325 ( .A1(n24436), .A2(n24435), .ZN(n24556) );
NAND2_X4 U34326 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n24554) );
OR2_X4 U34327 ( .A1(n24556), .A2(n20264), .ZN(n24438) );
NAND2_X4 U34328 ( .A1(n20264), .A2(n24556), .ZN(n24437) );
NAND2_X4 U34329 ( .A1(n24438), .A2(n24437), .ZN(n24493) );
NAND2_X4 U34330 ( .A1(n20340), .A2(n24439), .ZN(n24444) );
NAND2_X4 U34331 ( .A1(n20376), .A2(n24440), .ZN(n24442) );
NAND2_X4 U34332 ( .A1(n24442), .A2(n24441), .ZN(n24443) );
NAND2_X4 U34333 ( .A1(n24444), .A2(n24443), .ZN(n24564) );
NAND2_X4 U34334 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n24563) );
OR2_X4 U34335 ( .A1(n24564), .A2(n20301), .ZN(n24446) );
NAND2_X4 U34336 ( .A1(n20301), .A2(n24564), .ZN(n24445) );
NAND2_X4 U34337 ( .A1(n24446), .A2(n24445), .ZN(n24490) );
NAND2_X4 U34338 ( .A1(n20377), .A2(n20413), .ZN(n24452) );
NAND2_X4 U34339 ( .A1(n24448), .A2(n24447), .ZN(n24450) );
NAND2_X4 U34340 ( .A1(n24450), .A2(n24449), .ZN(n24451) );
NAND2_X4 U34341 ( .A1(n24452), .A2(n24451), .ZN(n24572) );
NAND2_X4 U34342 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n24570) );
OR2_X4 U34343 ( .A1(n24572), .A2(n20338), .ZN(n24454) );
NAND2_X4 U34344 ( .A1(n20338), .A2(n24572), .ZN(n24453) );
NAND2_X4 U34345 ( .A1(n24454), .A2(n24453), .ZN(n24487) );
NAND2_X4 U34346 ( .A1(n20414), .A2(n24455), .ZN(n24460) );
NAND2_X4 U34347 ( .A1(n20451), .A2(n24456), .ZN(n24458) );
NAND2_X4 U34348 ( .A1(n24458), .A2(n24457), .ZN(n24459) );
NAND2_X4 U34349 ( .A1(n24460), .A2(n24459), .ZN(n24580) );
NAND2_X4 U34350 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n24579) );
OR2_X4 U34351 ( .A1(n24580), .A2(n20375), .ZN(n24462) );
NAND2_X4 U34352 ( .A1(n20375), .A2(n24580), .ZN(n24461) );
NAND2_X4 U34353 ( .A1(n24462), .A2(n24461), .ZN(n24484) );
NAND2_X4 U34354 ( .A1(n20452), .A2(n20489), .ZN(n24468) );
NAND2_X4 U34355 ( .A1(n24464), .A2(n24463), .ZN(n24466) );
NAND2_X4 U34356 ( .A1(n24466), .A2(n24465), .ZN(n24467) );
NAND2_X4 U34357 ( .A1(n24468), .A2(n24467), .ZN(n24588) );
NAND2_X4 U34358 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n24586) );
OR2_X4 U34359 ( .A1(n24588), .A2(n20412), .ZN(n24470) );
NAND2_X4 U34360 ( .A1(n20412), .A2(n24588), .ZN(n24469) );
NAND2_X4 U34361 ( .A1(n24470), .A2(n24469), .ZN(n24481) );
NOR2_X4 U34362 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_5), .ZN(n24597) );
NAND2_X4 U34363 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n24596) );
NAND2_X4 U34364 ( .A1(n24597), .A2(n24596), .ZN(n24472) );
OR2_X4 U34365 ( .A1(n24596), .A2(n24597), .ZN(n24471) );
NAND2_X4 U34366 ( .A1(n24472), .A2(n24471), .ZN(n24478) );
NAND2_X4 U34367 ( .A1(n24474), .A2(n20490), .ZN(n24477) );
NAND2_X4 U34368 ( .A1(n20490), .A2(n24475), .ZN(n24476) );
NAND2_X4 U34369 ( .A1(n24477), .A2(n24476), .ZN(n24598) );
NAND2_X4 U34370 ( .A1(n24478), .A2(n24598), .ZN(n24480) );
OR2_X4 U34371 ( .A1(n24598), .A2(n24478), .ZN(n24479) );
NAND2_X4 U34372 ( .A1(n24480), .A2(n24479), .ZN(n24587) );
NAND2_X4 U34373 ( .A1(n24481), .A2(n20449), .ZN(n24483) );
OR2_X4 U34374 ( .A1(n20449), .A2(n24481), .ZN(n24482) );
NAND2_X4 U34375 ( .A1(n24483), .A2(n24482), .ZN(n24578) );
NAND2_X4 U34376 ( .A1(n24484), .A2(n20411), .ZN(n24486) );
OR2_X4 U34377 ( .A1(n20411), .A2(n24484), .ZN(n24485) );
NAND2_X4 U34378 ( .A1(n24486), .A2(n24485), .ZN(n24571) );
NAND2_X4 U34379 ( .A1(n24487), .A2(n20374), .ZN(n24489) );
OR2_X4 U34380 ( .A1(n20374), .A2(n24487), .ZN(n24488) );
NAND2_X4 U34381 ( .A1(n24489), .A2(n24488), .ZN(n24562) );
NAND2_X4 U34382 ( .A1(n24490), .A2(n20337), .ZN(n24492) );
OR2_X4 U34383 ( .A1(n20337), .A2(n24490), .ZN(n24491) );
NAND2_X4 U34384 ( .A1(n24492), .A2(n24491), .ZN(n24555) );
NAND2_X4 U34385 ( .A1(n24493), .A2(n20300), .ZN(n24495) );
OR2_X4 U34386 ( .A1(n20300), .A2(n24493), .ZN(n24494) );
NAND2_X4 U34387 ( .A1(n24495), .A2(n24494), .ZN(n24546) );
NAND2_X4 U34388 ( .A1(n24496), .A2(n20263), .ZN(n24498) );
OR2_X4 U34389 ( .A1(n20263), .A2(n24496), .ZN(n24497) );
NAND2_X4 U34390 ( .A1(n24498), .A2(n24497), .ZN(n24539) );
NAND2_X4 U34391 ( .A1(n24499), .A2(n20227), .ZN(n24501) );
OR2_X4 U34392 ( .A1(n20227), .A2(n24499), .ZN(n24500) );
NAND2_X4 U34393 ( .A1(n24501), .A2(n24500), .ZN(n24530) );
NAND2_X4 U34394 ( .A1(n24502), .A2(n20191), .ZN(n24504) );
OR2_X4 U34395 ( .A1(n20191), .A2(n24502), .ZN(n24503) );
NAND2_X4 U34396 ( .A1(n24504), .A2(n24503), .ZN(n24629) );
NAND2_X4 U34397 ( .A1(n24505), .A2(n20155), .ZN(n24507) );
OR2_X4 U34398 ( .A1(n20155), .A2(n24505), .ZN(n24506) );
NAND2_X4 U34399 ( .A1(n24507), .A2(n24506), .ZN(n24639) );
NAND2_X4 U34400 ( .A1(n20101), .A2(n24508), .ZN(n24513) );
NAND2_X4 U34401 ( .A1(n20157), .A2(n24509), .ZN(n24511) );
NAND2_X4 U34402 ( .A1(n24511), .A2(n24510), .ZN(n24512) );
NAND2_X4 U34403 ( .A1(n24513), .A2(n24512), .ZN(n24638) );
NOR2_X4 U34404 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_5), .ZN(n24637) );
NOR2_X4 U34405 ( .A1(n24638), .A2(n24637), .ZN(n24514) );
OR2_X4 U34406 ( .A1(n20099), .A2(n24514), .ZN(n24516) );
NAND2_X4 U34407 ( .A1(n24514), .A2(n20099), .ZN(n24515) );
NAND2_X4 U34408 ( .A1(n24516), .A2(n24515), .ZN(n25248) );
NAND2_X4 U34409 ( .A1(n24517), .A2(n24519), .ZN(n24521) );
NAND2_X4 U34410 ( .A1(n24519), .A2(n24518), .ZN(n24520) );
NAND2_X4 U34411 ( .A1(n24521), .A2(n24520), .ZN(n25247) );
NAND2_X4 U34412 ( .A1(n25248), .A2(n25247), .ZN(n24523) );
OR2_X4 U34413 ( .A1(n25247), .A2(n25248), .ZN(n24522) );
NAND2_X4 U34414 ( .A1(n24523), .A2(n24522), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_19_) );
OR2_X4 U34415 ( .A1(n24524), .A2(n20586), .ZN(n24526) );
NAND2_X4 U34416 ( .A1(n20586), .A2(n24524), .ZN(n24525) );
NAND2_X4 U34417 ( .A1(n24526), .A2(n24525), .ZN(n24527) );
NOR2_X4 U34418 ( .A1(n24527), .A2(n20622), .ZN(n24529) );
AND2_X4 U34419 ( .A1(n20622), .A2(n24527), .ZN(n24528) );
NOR2_X4 U34420 ( .A1(n24529), .A2(n24528), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N38) );
NAND2_X4 U34421 ( .A1(n20156), .A2(n24530), .ZN(n24535) );
NAND2_X4 U34422 ( .A1(n20191), .A2(n24531), .ZN(n24533) );
NAND2_X4 U34423 ( .A1(n24533), .A2(n24532), .ZN(n24534) );
NAND2_X4 U34424 ( .A1(n24535), .A2(n24534), .ZN(n24734) );
NAND2_X4 U34425 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n24733) );
OR2_X4 U34426 ( .A1(n24734), .A2(n20098), .ZN(n24537) );
NAND2_X4 U34427 ( .A1(n20098), .A2(n24734), .ZN(n24536) );
NAND2_X4 U34428 ( .A1(n24537), .A2(n24536), .ZN(n24625) );
NAND2_X4 U34429 ( .A1(n20192), .A2(n20227), .ZN(n24543) );
NAND2_X4 U34430 ( .A1(n24539), .A2(n24538), .ZN(n24541) );
NAND2_X4 U34431 ( .A1(n24541), .A2(n24540), .ZN(n24542) );
NAND2_X4 U34432 ( .A1(n24543), .A2(n24542), .ZN(n24647) );
NAND2_X4 U34433 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n24645) );
OR2_X4 U34434 ( .A1(n24647), .A2(n20154), .ZN(n24545) );
NAND2_X4 U34435 ( .A1(n20154), .A2(n24647), .ZN(n24544) );
NAND2_X4 U34436 ( .A1(n24545), .A2(n24544), .ZN(n24622) );
NAND2_X4 U34437 ( .A1(n20228), .A2(n24546), .ZN(n24551) );
NAND2_X4 U34438 ( .A1(n20263), .A2(n24547), .ZN(n24549) );
NAND2_X4 U34439 ( .A1(n24549), .A2(n24548), .ZN(n24550) );
NAND2_X4 U34440 ( .A1(n24551), .A2(n24550), .ZN(n24655) );
NAND2_X4 U34441 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n24654) );
OR2_X4 U34442 ( .A1(n24655), .A2(n20190), .ZN(n24553) );
NAND2_X4 U34443 ( .A1(n20190), .A2(n24655), .ZN(n24552) );
NAND2_X4 U34444 ( .A1(n24553), .A2(n24552), .ZN(n24619) );
NAND2_X4 U34445 ( .A1(n20264), .A2(n20300), .ZN(n24559) );
NAND2_X4 U34446 ( .A1(n24555), .A2(n24554), .ZN(n24557) );
NAND2_X4 U34447 ( .A1(n24557), .A2(n24556), .ZN(n24558) );
NAND2_X4 U34448 ( .A1(n24559), .A2(n24558), .ZN(n24663) );
NAND2_X4 U34449 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n24661) );
OR2_X4 U34450 ( .A1(n24663), .A2(n20226), .ZN(n24561) );
NAND2_X4 U34451 ( .A1(n20226), .A2(n24663), .ZN(n24560) );
NAND2_X4 U34452 ( .A1(n24561), .A2(n24560), .ZN(n24616) );
NAND2_X4 U34453 ( .A1(n20301), .A2(n24562), .ZN(n24567) );
NAND2_X4 U34454 ( .A1(n20337), .A2(n24563), .ZN(n24565) );
NAND2_X4 U34455 ( .A1(n24565), .A2(n24564), .ZN(n24566) );
NAND2_X4 U34456 ( .A1(n24567), .A2(n24566), .ZN(n24671) );
NAND2_X4 U34457 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n24670) );
OR2_X4 U34458 ( .A1(n24671), .A2(n20262), .ZN(n24569) );
NAND2_X4 U34459 ( .A1(n20262), .A2(n24671), .ZN(n24568) );
NAND2_X4 U34460 ( .A1(n24569), .A2(n24568), .ZN(n24613) );
NAND2_X4 U34461 ( .A1(n20338), .A2(n20374), .ZN(n24575) );
NAND2_X4 U34462 ( .A1(n24571), .A2(n24570), .ZN(n24573) );
NAND2_X4 U34463 ( .A1(n24573), .A2(n24572), .ZN(n24574) );
NAND2_X4 U34464 ( .A1(n24575), .A2(n24574), .ZN(n24679) );
NAND2_X4 U34465 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n24677) );
OR2_X4 U34466 ( .A1(n24679), .A2(n20299), .ZN(n24577) );
NAND2_X4 U34467 ( .A1(n20299), .A2(n24679), .ZN(n24576) );
NAND2_X4 U34468 ( .A1(n24577), .A2(n24576), .ZN(n24610) );
NAND2_X4 U34469 ( .A1(n20375), .A2(n24578), .ZN(n24583) );
NAND2_X4 U34470 ( .A1(n20411), .A2(n24579), .ZN(n24581) );
NAND2_X4 U34471 ( .A1(n24581), .A2(n24580), .ZN(n24582) );
NAND2_X4 U34472 ( .A1(n24583), .A2(n24582), .ZN(n24687) );
NAND2_X4 U34473 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n24686) );
OR2_X4 U34474 ( .A1(n24687), .A2(n20336), .ZN(n24585) );
NAND2_X4 U34475 ( .A1(n20336), .A2(n24687), .ZN(n24584) );
NAND2_X4 U34476 ( .A1(n24585), .A2(n24584), .ZN(n24607) );
NAND2_X4 U34477 ( .A1(n20412), .A2(n20449), .ZN(n24591) );
NAND2_X4 U34478 ( .A1(n24587), .A2(n24586), .ZN(n24589) );
NAND2_X4 U34479 ( .A1(n24589), .A2(n24588), .ZN(n24590) );
NAND2_X4 U34480 ( .A1(n24591), .A2(n24590), .ZN(n24695) );
NAND2_X4 U34481 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n24693) );
OR2_X4 U34482 ( .A1(n24695), .A2(n20373), .ZN(n24593) );
NAND2_X4 U34483 ( .A1(n20373), .A2(n24695), .ZN(n24592) );
NAND2_X4 U34484 ( .A1(n24593), .A2(n24592), .ZN(n24604) );
NOR2_X4 U34485 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_6), .ZN(n24704) );
NAND2_X4 U34486 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n24703) );
NAND2_X4 U34487 ( .A1(n24704), .A2(n24703), .ZN(n24595) );
OR2_X4 U34488 ( .A1(n24703), .A2(n24704), .ZN(n24594) );
NAND2_X4 U34489 ( .A1(n24595), .A2(n24594), .ZN(n24601) );
NAND2_X4 U34490 ( .A1(n24597), .A2(n20450), .ZN(n24600) );
NAND2_X4 U34491 ( .A1(n20450), .A2(n24598), .ZN(n24599) );
NAND2_X4 U34492 ( .A1(n24600), .A2(n24599), .ZN(n24705) );
NAND2_X4 U34493 ( .A1(n24601), .A2(n24705), .ZN(n24603) );
OR2_X4 U34494 ( .A1(n24705), .A2(n24601), .ZN(n24602) );
NAND2_X4 U34495 ( .A1(n24603), .A2(n24602), .ZN(n24694) );
NAND2_X4 U34496 ( .A1(n24604), .A2(n20409), .ZN(n24606) );
OR2_X4 U34497 ( .A1(n20409), .A2(n24604), .ZN(n24605) );
NAND2_X4 U34498 ( .A1(n24606), .A2(n24605), .ZN(n24685) );
NAND2_X4 U34499 ( .A1(n24607), .A2(n20372), .ZN(n24609) );
OR2_X4 U34500 ( .A1(n20372), .A2(n24607), .ZN(n24608) );
NAND2_X4 U34501 ( .A1(n24609), .A2(n24608), .ZN(n24678) );
NAND2_X4 U34502 ( .A1(n24610), .A2(n20335), .ZN(n24612) );
OR2_X4 U34503 ( .A1(n20335), .A2(n24610), .ZN(n24611) );
NAND2_X4 U34504 ( .A1(n24612), .A2(n24611), .ZN(n24669) );
NAND2_X4 U34505 ( .A1(n24613), .A2(n20298), .ZN(n24615) );
OR2_X4 U34506 ( .A1(n20298), .A2(n24613), .ZN(n24614) );
NAND2_X4 U34507 ( .A1(n24615), .A2(n24614), .ZN(n24662) );
NAND2_X4 U34508 ( .A1(n24616), .A2(n20261), .ZN(n24618) );
OR2_X4 U34509 ( .A1(n20261), .A2(n24616), .ZN(n24617) );
NAND2_X4 U34510 ( .A1(n24618), .A2(n24617), .ZN(n24653) );
NAND2_X4 U34511 ( .A1(n24619), .A2(n20225), .ZN(n24621) );
OR2_X4 U34512 ( .A1(n20225), .A2(n24619), .ZN(n24620) );
NAND2_X4 U34513 ( .A1(n24621), .A2(n24620), .ZN(n24646) );
NAND2_X4 U34514 ( .A1(n24622), .A2(n20189), .ZN(n24624) );
OR2_X4 U34515 ( .A1(n20189), .A2(n24622), .ZN(n24623) );
NAND2_X4 U34516 ( .A1(n24624), .A2(n24623), .ZN(n24732) );
NAND2_X4 U34517 ( .A1(n24625), .A2(n20153), .ZN(n24627) );
OR2_X4 U34518 ( .A1(n20153), .A2(n24625), .ZN(n24626) );
AND2_X4 U34519 ( .A1(n24627), .A2(n24626), .ZN(n24743) );
NAND2_X4 U34520 ( .A1(n20100), .A2(n20155), .ZN(n24633) );
NAND2_X4 U34521 ( .A1(n24629), .A2(n24628), .ZN(n24631) );
NAND2_X4 U34522 ( .A1(n24631), .A2(n24630), .ZN(n24632) );
NAND2_X4 U34523 ( .A1(n24633), .A2(n24632), .ZN(n24742) );
NOR2_X4 U34524 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_6), .ZN(n24741) );
NOR2_X4 U34525 ( .A1(n24742), .A2(n24741), .ZN(n24634) );
OR2_X4 U34526 ( .A1(n24743), .A2(n24634), .ZN(n24636) );
NAND2_X4 U34527 ( .A1(n24634), .A2(n24743), .ZN(n24635) );
NAND2_X4 U34528 ( .A1(n24636), .A2(n24635), .ZN(n24643) );
NAND2_X4 U34529 ( .A1(n24637), .A2(n24639), .ZN(n24641) );
NAND2_X4 U34530 ( .A1(n24639), .A2(n24638), .ZN(n24640) );
NAND2_X4 U34531 ( .A1(n24641), .A2(n24640), .ZN(n24642) );
NOR2_X4 U34532 ( .A1(n24643), .A2(n24642), .ZN(n24644) );
NOR2_X4 U34533 ( .A1(n20063), .A2(n20062), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_21_) );
NOR2_X4 U34534 ( .A1(n24644), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_21_), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_20_) );
NAND2_X4 U34535 ( .A1(n20154), .A2(n20189), .ZN(n24650) );
NAND2_X4 U34536 ( .A1(n24646), .A2(n24645), .ZN(n24648) );
NAND2_X4 U34537 ( .A1(n24648), .A2(n24647), .ZN(n24649) );
NAND2_X4 U34538 ( .A1(n24650), .A2(n24649), .ZN(n24826) );
NAND2_X4 U34539 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n24824) );
OR2_X4 U34540 ( .A1(n24826), .A2(n20097), .ZN(n24652) );
NAND2_X4 U34541 ( .A1(n20097), .A2(n24826), .ZN(n24651) );
NAND2_X4 U34542 ( .A1(n24652), .A2(n24651), .ZN(n24729) );
NAND2_X4 U34543 ( .A1(n20190), .A2(n24653), .ZN(n24658) );
NAND2_X4 U34544 ( .A1(n20225), .A2(n24654), .ZN(n24656) );
NAND2_X4 U34545 ( .A1(n24656), .A2(n24655), .ZN(n24657) );
NAND2_X4 U34546 ( .A1(n24658), .A2(n24657), .ZN(n24750) );
NAND2_X4 U34547 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n24749) );
OR2_X4 U34548 ( .A1(n24750), .A2(n20152), .ZN(n24660) );
NAND2_X4 U34549 ( .A1(n20152), .A2(n24750), .ZN(n24659) );
NAND2_X4 U34550 ( .A1(n24660), .A2(n24659), .ZN(n24726) );
NAND2_X4 U34551 ( .A1(n20226), .A2(n20261), .ZN(n24666) );
NAND2_X4 U34552 ( .A1(n24662), .A2(n24661), .ZN(n24664) );
NAND2_X4 U34553 ( .A1(n24664), .A2(n24663), .ZN(n24665) );
NAND2_X4 U34554 ( .A1(n24666), .A2(n24665), .ZN(n24758) );
NAND2_X4 U34555 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n24756) );
OR2_X4 U34556 ( .A1(n24758), .A2(n20188), .ZN(n24668) );
NAND2_X4 U34557 ( .A1(n20188), .A2(n24758), .ZN(n24667) );
NAND2_X4 U34558 ( .A1(n24668), .A2(n24667), .ZN(n24723) );
NAND2_X4 U34559 ( .A1(n20262), .A2(n24669), .ZN(n24674) );
NAND2_X4 U34560 ( .A1(n20298), .A2(n24670), .ZN(n24672) );
NAND2_X4 U34561 ( .A1(n24672), .A2(n24671), .ZN(n24673) );
NAND2_X4 U34562 ( .A1(n24674), .A2(n24673), .ZN(n24766) );
NAND2_X4 U34563 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n24765) );
OR2_X4 U34564 ( .A1(n24766), .A2(n20224), .ZN(n24676) );
NAND2_X4 U34565 ( .A1(n20224), .A2(n24766), .ZN(n24675) );
NAND2_X4 U34566 ( .A1(n24676), .A2(n24675), .ZN(n24720) );
NAND2_X4 U34567 ( .A1(n20299), .A2(n20335), .ZN(n24682) );
NAND2_X4 U34568 ( .A1(n24678), .A2(n24677), .ZN(n24680) );
NAND2_X4 U34569 ( .A1(n24680), .A2(n24679), .ZN(n24681) );
NAND2_X4 U34570 ( .A1(n24682), .A2(n24681), .ZN(n24774) );
NAND2_X4 U34571 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n24772) );
OR2_X4 U34572 ( .A1(n24774), .A2(n20260), .ZN(n24684) );
NAND2_X4 U34573 ( .A1(n20260), .A2(n24774), .ZN(n24683) );
NAND2_X4 U34574 ( .A1(n24684), .A2(n24683), .ZN(n24717) );
NAND2_X4 U34575 ( .A1(n20336), .A2(n24685), .ZN(n24690) );
NAND2_X4 U34576 ( .A1(n20372), .A2(n24686), .ZN(n24688) );
NAND2_X4 U34577 ( .A1(n24688), .A2(n24687), .ZN(n24689) );
NAND2_X4 U34578 ( .A1(n24690), .A2(n24689), .ZN(n24782) );
NAND2_X4 U34579 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n24781) );
OR2_X4 U34580 ( .A1(n24782), .A2(n20297), .ZN(n24692) );
NAND2_X4 U34581 ( .A1(n20297), .A2(n24782), .ZN(n24691) );
NAND2_X4 U34582 ( .A1(n24692), .A2(n24691), .ZN(n24714) );
NAND2_X4 U34583 ( .A1(n20373), .A2(n20409), .ZN(n24698) );
NAND2_X4 U34584 ( .A1(n24694), .A2(n24693), .ZN(n24696) );
NAND2_X4 U34585 ( .A1(n24696), .A2(n24695), .ZN(n24697) );
NAND2_X4 U34586 ( .A1(n24698), .A2(n24697), .ZN(n24790) );
NAND2_X4 U34587 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n24788) );
OR2_X4 U34588 ( .A1(n24790), .A2(n20334), .ZN(n24700) );
NAND2_X4 U34589 ( .A1(n20334), .A2(n24790), .ZN(n24699) );
NAND2_X4 U34590 ( .A1(n24700), .A2(n24699), .ZN(n24711) );
NOR2_X4 U34591 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_7), .ZN(n24799) );
NAND2_X4 U34592 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n24798) );
NAND2_X4 U34593 ( .A1(n24799), .A2(n24798), .ZN(n24702) );
OR2_X4 U34594 ( .A1(n24798), .A2(n24799), .ZN(n24701) );
NAND2_X4 U34595 ( .A1(n24702), .A2(n24701), .ZN(n24708) );
NAND2_X4 U34596 ( .A1(n24704), .A2(n20410), .ZN(n24707) );
NAND2_X4 U34597 ( .A1(n20410), .A2(n24705), .ZN(n24706) );
NAND2_X4 U34598 ( .A1(n24707), .A2(n24706), .ZN(n24800) );
NAND2_X4 U34599 ( .A1(n24708), .A2(n24800), .ZN(n24710) );
OR2_X4 U34600 ( .A1(n24800), .A2(n24708), .ZN(n24709) );
NAND2_X4 U34601 ( .A1(n24710), .A2(n24709), .ZN(n24789) );
NAND2_X4 U34602 ( .A1(n24711), .A2(n20370), .ZN(n24713) );
OR2_X4 U34603 ( .A1(n20370), .A2(n24711), .ZN(n24712) );
NAND2_X4 U34604 ( .A1(n24713), .A2(n24712), .ZN(n24780) );
NAND2_X4 U34605 ( .A1(n24714), .A2(n20333), .ZN(n24716) );
OR2_X4 U34606 ( .A1(n20333), .A2(n24714), .ZN(n24715) );
NAND2_X4 U34607 ( .A1(n24716), .A2(n24715), .ZN(n24773) );
NAND2_X4 U34608 ( .A1(n24717), .A2(n20296), .ZN(n24719) );
OR2_X4 U34609 ( .A1(n20296), .A2(n24717), .ZN(n24718) );
NAND2_X4 U34610 ( .A1(n24719), .A2(n24718), .ZN(n24764) );
NAND2_X4 U34611 ( .A1(n24720), .A2(n20259), .ZN(n24722) );
OR2_X4 U34612 ( .A1(n20259), .A2(n24720), .ZN(n24721) );
NAND2_X4 U34613 ( .A1(n24722), .A2(n24721), .ZN(n24757) );
NAND2_X4 U34614 ( .A1(n24723), .A2(n20223), .ZN(n24725) );
OR2_X4 U34615 ( .A1(n20223), .A2(n24723), .ZN(n24724) );
NAND2_X4 U34616 ( .A1(n24725), .A2(n24724), .ZN(n24748) );
NAND2_X4 U34617 ( .A1(n24726), .A2(n20187), .ZN(n24728) );
OR2_X4 U34618 ( .A1(n20187), .A2(n24726), .ZN(n24727) );
NAND2_X4 U34619 ( .A1(n24728), .A2(n24727), .ZN(n24825) );
NAND2_X4 U34620 ( .A1(n24729), .A2(n20151), .ZN(n24731) );
OR2_X4 U34621 ( .A1(n20151), .A2(n24729), .ZN(n24730) );
NAND2_X4 U34622 ( .A1(n24731), .A2(n24730), .ZN(n24835) );
NAND2_X4 U34623 ( .A1(n20098), .A2(n24732), .ZN(n24737) );
NAND2_X4 U34624 ( .A1(n20153), .A2(n24733), .ZN(n24735) );
NAND2_X4 U34625 ( .A1(n24735), .A2(n24734), .ZN(n24736) );
NAND2_X4 U34626 ( .A1(n24737), .A2(n24736), .ZN(n24834) );
NOR2_X4 U34627 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_7), .ZN(n24833) );
NOR2_X4 U34628 ( .A1(n24834), .A2(n24833), .ZN(n24738) );
OR2_X4 U34629 ( .A1(n20096), .A2(n24738), .ZN(n24740) );
NAND2_X4 U34630 ( .A1(n24738), .A2(n20096), .ZN(n24739) );
NAND2_X4 U34631 ( .A1(n24740), .A2(n24739), .ZN(n25250) );
NAND2_X4 U34632 ( .A1(n24741), .A2(n24743), .ZN(n24745) );
NAND2_X4 U34633 ( .A1(n24743), .A2(n24742), .ZN(n24744) );
NAND2_X4 U34634 ( .A1(n24745), .A2(n24744), .ZN(n25249) );
NAND2_X4 U34635 ( .A1(n25250), .A2(n25249), .ZN(n24747) );
OR2_X4 U34636 ( .A1(n25249), .A2(n25250), .ZN(n24746) );
NAND2_X4 U34637 ( .A1(n24747), .A2(n24746), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_21_) );
NAND2_X4 U34638 ( .A1(n20152), .A2(n24748), .ZN(n24753) );
NAND2_X4 U34639 ( .A1(n20187), .A2(n24749), .ZN(n24751) );
NAND2_X4 U34640 ( .A1(n24751), .A2(n24750), .ZN(n24752) );
NAND2_X4 U34641 ( .A1(n24753), .A2(n24752), .ZN(n24908) );
NAND2_X4 U34642 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n24907) );
OR2_X4 U34643 ( .A1(n24908), .A2(n20095), .ZN(n24755) );
NAND2_X4 U34644 ( .A1(n20095), .A2(n24908), .ZN(n24754) );
NAND2_X4 U34645 ( .A1(n24755), .A2(n24754), .ZN(n24821) );
NAND2_X4 U34646 ( .A1(n20188), .A2(n20223), .ZN(n24761) );
NAND2_X4 U34647 ( .A1(n24757), .A2(n24756), .ZN(n24759) );
NAND2_X4 U34648 ( .A1(n24759), .A2(n24758), .ZN(n24760) );
NAND2_X4 U34649 ( .A1(n24761), .A2(n24760), .ZN(n24843) );
NAND2_X4 U34650 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n24841) );
OR2_X4 U34651 ( .A1(n24843), .A2(n20150), .ZN(n24763) );
NAND2_X4 U34652 ( .A1(n20150), .A2(n24843), .ZN(n24762) );
NAND2_X4 U34653 ( .A1(n24763), .A2(n24762), .ZN(n24818) );
NAND2_X4 U34654 ( .A1(n20224), .A2(n24764), .ZN(n24769) );
NAND2_X4 U34655 ( .A1(n20259), .A2(n24765), .ZN(n24767) );
NAND2_X4 U34656 ( .A1(n24767), .A2(n24766), .ZN(n24768) );
NAND2_X4 U34657 ( .A1(n24769), .A2(n24768), .ZN(n24851) );
NAND2_X4 U34658 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n24850) );
OR2_X4 U34659 ( .A1(n24851), .A2(n20186), .ZN(n24771) );
NAND2_X4 U34660 ( .A1(n20186), .A2(n24851), .ZN(n24770) );
NAND2_X4 U34661 ( .A1(n24771), .A2(n24770), .ZN(n24815) );
NAND2_X4 U34662 ( .A1(n20260), .A2(n20296), .ZN(n24777) );
NAND2_X4 U34663 ( .A1(n24773), .A2(n24772), .ZN(n24775) );
NAND2_X4 U34664 ( .A1(n24775), .A2(n24774), .ZN(n24776) );
NAND2_X4 U34665 ( .A1(n24777), .A2(n24776), .ZN(n24859) );
NAND2_X4 U34666 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n24857) );
OR2_X4 U34667 ( .A1(n24859), .A2(n20222), .ZN(n24779) );
NAND2_X4 U34668 ( .A1(n20222), .A2(n24859), .ZN(n24778) );
NAND2_X4 U34669 ( .A1(n24779), .A2(n24778), .ZN(n24812) );
NAND2_X4 U34670 ( .A1(n20297), .A2(n24780), .ZN(n24785) );
NAND2_X4 U34671 ( .A1(n20333), .A2(n24781), .ZN(n24783) );
NAND2_X4 U34672 ( .A1(n24783), .A2(n24782), .ZN(n24784) );
NAND2_X4 U34673 ( .A1(n24785), .A2(n24784), .ZN(n24867) );
NAND2_X4 U34674 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n24866) );
OR2_X4 U34675 ( .A1(n24867), .A2(n20258), .ZN(n24787) );
NAND2_X4 U34676 ( .A1(n20258), .A2(n24867), .ZN(n24786) );
NAND2_X4 U34677 ( .A1(n24787), .A2(n24786), .ZN(n24809) );
NAND2_X4 U34678 ( .A1(n20334), .A2(n20370), .ZN(n24793) );
NAND2_X4 U34679 ( .A1(n24789), .A2(n24788), .ZN(n24791) );
NAND2_X4 U34680 ( .A1(n24791), .A2(n24790), .ZN(n24792) );
NAND2_X4 U34681 ( .A1(n24793), .A2(n24792), .ZN(n24875) );
NAND2_X4 U34682 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n24873) );
OR2_X4 U34683 ( .A1(n24875), .A2(n20295), .ZN(n24795) );
NAND2_X4 U34684 ( .A1(n20295), .A2(n24875), .ZN(n24794) );
NAND2_X4 U34685 ( .A1(n24795), .A2(n24794), .ZN(n24806) );
NOR2_X4 U34686 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_8), .ZN(n24884) );
NAND2_X4 U34687 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n24883) );
NAND2_X4 U34688 ( .A1(n24884), .A2(n24883), .ZN(n24797) );
OR2_X4 U34689 ( .A1(n24883), .A2(n24884), .ZN(n24796) );
NAND2_X4 U34690 ( .A1(n24797), .A2(n24796), .ZN(n24803) );
NAND2_X4 U34691 ( .A1(n24799), .A2(n20371), .ZN(n24802) );
NAND2_X4 U34692 ( .A1(n20371), .A2(n24800), .ZN(n24801) );
NAND2_X4 U34693 ( .A1(n24802), .A2(n24801), .ZN(n24885) );
NAND2_X4 U34694 ( .A1(n24803), .A2(n24885), .ZN(n24805) );
OR2_X4 U34695 ( .A1(n24885), .A2(n24803), .ZN(n24804) );
NAND2_X4 U34696 ( .A1(n24805), .A2(n24804), .ZN(n24874) );
NAND2_X4 U34697 ( .A1(n24806), .A2(n20331), .ZN(n24808) );
OR2_X4 U34698 ( .A1(n20331), .A2(n24806), .ZN(n24807) );
NAND2_X4 U34699 ( .A1(n24808), .A2(n24807), .ZN(n24865) );
NAND2_X4 U34700 ( .A1(n24809), .A2(n20294), .ZN(n24811) );
OR2_X4 U34701 ( .A1(n20294), .A2(n24809), .ZN(n24810) );
NAND2_X4 U34702 ( .A1(n24811), .A2(n24810), .ZN(n24858) );
NAND2_X4 U34703 ( .A1(n24812), .A2(n20257), .ZN(n24814) );
OR2_X4 U34704 ( .A1(n20257), .A2(n24812), .ZN(n24813) );
NAND2_X4 U34705 ( .A1(n24814), .A2(n24813), .ZN(n24849) );
NAND2_X4 U34706 ( .A1(n24815), .A2(n20221), .ZN(n24817) );
OR2_X4 U34707 ( .A1(n20221), .A2(n24815), .ZN(n24816) );
NAND2_X4 U34708 ( .A1(n24817), .A2(n24816), .ZN(n24842) );
NAND2_X4 U34709 ( .A1(n24818), .A2(n20185), .ZN(n24820) );
OR2_X4 U34710 ( .A1(n20185), .A2(n24818), .ZN(n24819) );
NAND2_X4 U34711 ( .A1(n24820), .A2(n24819), .ZN(n24906) );
NAND2_X4 U34712 ( .A1(n24821), .A2(n20149), .ZN(n24823) );
OR2_X4 U34713 ( .A1(n20149), .A2(n24821), .ZN(n24822) );
AND2_X4 U34714 ( .A1(n24823), .A2(n24822), .ZN(n24917) );
NAND2_X4 U34715 ( .A1(n20097), .A2(n20151), .ZN(n24829) );
NAND2_X4 U34716 ( .A1(n24825), .A2(n24824), .ZN(n24827) );
NAND2_X4 U34717 ( .A1(n24827), .A2(n24826), .ZN(n24828) );
NAND2_X4 U34718 ( .A1(n24829), .A2(n24828), .ZN(n24916) );
NOR2_X4 U34719 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_8), .ZN(n24915) );
NOR2_X4 U34720 ( .A1(n24916), .A2(n24915), .ZN(n24830) );
OR2_X4 U34721 ( .A1(n24917), .A2(n24830), .ZN(n24832) );
NAND2_X4 U34722 ( .A1(n24830), .A2(n24917), .ZN(n24831) );
NAND2_X4 U34723 ( .A1(n24832), .A2(n24831), .ZN(n24839) );
NAND2_X4 U34724 ( .A1(n24833), .A2(n24835), .ZN(n24837) );
NAND2_X4 U34725 ( .A1(n24835), .A2(n24834), .ZN(n24836) );
NAND2_X4 U34726 ( .A1(n24837), .A2(n24836), .ZN(n24838) );
NOR2_X4 U34727 ( .A1(n24839), .A2(n24838), .ZN(n24840) );
NOR2_X4 U34728 ( .A1(n20056), .A2(n20055), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_23_) );
NOR2_X4 U34729 ( .A1(n24840), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_23_), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_22_) );
NAND2_X4 U34730 ( .A1(n20150), .A2(n20185), .ZN(n24846) );
NAND2_X4 U34731 ( .A1(n24842), .A2(n24841), .ZN(n24844) );
NAND2_X4 U34732 ( .A1(n24844), .A2(n24843), .ZN(n24845) );
NAND2_X4 U34733 ( .A1(n24846), .A2(n24845), .ZN(n24978) );
NAND2_X4 U34734 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n24976) );
OR2_X4 U34735 ( .A1(n24978), .A2(n20094), .ZN(n24848) );
NAND2_X4 U34736 ( .A1(n20094), .A2(n24978), .ZN(n24847) );
NAND2_X4 U34737 ( .A1(n24848), .A2(n24847), .ZN(n24903) );
NAND2_X4 U34738 ( .A1(n20186), .A2(n24849), .ZN(n24854) );
NAND2_X4 U34739 ( .A1(n20221), .A2(n24850), .ZN(n24852) );
NAND2_X4 U34740 ( .A1(n24852), .A2(n24851), .ZN(n24853) );
NAND2_X4 U34741 ( .A1(n24854), .A2(n24853), .ZN(n24924) );
NAND2_X4 U34742 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n24923) );
OR2_X4 U34743 ( .A1(n24924), .A2(n20148), .ZN(n24856) );
NAND2_X4 U34744 ( .A1(n20148), .A2(n24924), .ZN(n24855) );
NAND2_X4 U34745 ( .A1(n24856), .A2(n24855), .ZN(n24900) );
NAND2_X4 U34746 ( .A1(n20222), .A2(n20257), .ZN(n24862) );
NAND2_X4 U34747 ( .A1(n24858), .A2(n24857), .ZN(n24860) );
NAND2_X4 U34748 ( .A1(n24860), .A2(n24859), .ZN(n24861) );
NAND2_X4 U34749 ( .A1(n24862), .A2(n24861), .ZN(n24932) );
NAND2_X4 U34750 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n24930) );
OR2_X4 U34751 ( .A1(n24932), .A2(n20184), .ZN(n24864) );
NAND2_X4 U34752 ( .A1(n20184), .A2(n24932), .ZN(n24863) );
NAND2_X4 U34753 ( .A1(n24864), .A2(n24863), .ZN(n24897) );
NAND2_X4 U34754 ( .A1(n20258), .A2(n24865), .ZN(n24870) );
NAND2_X4 U34755 ( .A1(n20294), .A2(n24866), .ZN(n24868) );
NAND2_X4 U34756 ( .A1(n24868), .A2(n24867), .ZN(n24869) );
NAND2_X4 U34757 ( .A1(n24870), .A2(n24869), .ZN(n24940) );
NAND2_X4 U34758 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n24939) );
OR2_X4 U34759 ( .A1(n24940), .A2(n20220), .ZN(n24872) );
NAND2_X4 U34760 ( .A1(n20220), .A2(n24940), .ZN(n24871) );
NAND2_X4 U34761 ( .A1(n24872), .A2(n24871), .ZN(n24894) );
NAND2_X4 U34762 ( .A1(n20295), .A2(n20331), .ZN(n24878) );
NAND2_X4 U34763 ( .A1(n24874), .A2(n24873), .ZN(n24876) );
NAND2_X4 U34764 ( .A1(n24876), .A2(n24875), .ZN(n24877) );
NAND2_X4 U34765 ( .A1(n24878), .A2(n24877), .ZN(n24948) );
NAND2_X4 U34766 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n24946) );
OR2_X4 U34767 ( .A1(n24948), .A2(n20256), .ZN(n24880) );
NAND2_X4 U34768 ( .A1(n20256), .A2(n24948), .ZN(n24879) );
NAND2_X4 U34769 ( .A1(n24880), .A2(n24879), .ZN(n24891) );
NOR2_X4 U34770 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_9), .ZN(n24957) );
NAND2_X4 U34771 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n24956) );
NAND2_X4 U34772 ( .A1(n24957), .A2(n24956), .ZN(n24882) );
OR2_X4 U34773 ( .A1(n24956), .A2(n24957), .ZN(n24881) );
NAND2_X4 U34774 ( .A1(n24882), .A2(n24881), .ZN(n24888) );
NAND2_X4 U34775 ( .A1(n24884), .A2(n20332), .ZN(n24887) );
NAND2_X4 U34776 ( .A1(n20332), .A2(n24885), .ZN(n24886) );
NAND2_X4 U34777 ( .A1(n24887), .A2(n24886), .ZN(n24958) );
NAND2_X4 U34778 ( .A1(n24888), .A2(n24958), .ZN(n24890) );
OR2_X4 U34779 ( .A1(n24958), .A2(n24888), .ZN(n24889) );
NAND2_X4 U34780 ( .A1(n24890), .A2(n24889), .ZN(n24947) );
NAND2_X4 U34781 ( .A1(n24891), .A2(n20292), .ZN(n24893) );
OR2_X4 U34782 ( .A1(n20292), .A2(n24891), .ZN(n24892) );
NAND2_X4 U34783 ( .A1(n24893), .A2(n24892), .ZN(n24938) );
NAND2_X4 U34784 ( .A1(n24894), .A2(n20255), .ZN(n24896) );
OR2_X4 U34785 ( .A1(n20255), .A2(n24894), .ZN(n24895) );
NAND2_X4 U34786 ( .A1(n24896), .A2(n24895), .ZN(n24931) );
NAND2_X4 U34787 ( .A1(n24897), .A2(n20219), .ZN(n24899) );
OR2_X4 U34788 ( .A1(n20219), .A2(n24897), .ZN(n24898) );
NAND2_X4 U34789 ( .A1(n24899), .A2(n24898), .ZN(n24922) );
NAND2_X4 U34790 ( .A1(n24900), .A2(n20183), .ZN(n24902) );
OR2_X4 U34791 ( .A1(n20183), .A2(n24900), .ZN(n24901) );
NAND2_X4 U34792 ( .A1(n24902), .A2(n24901), .ZN(n24977) );
NAND2_X4 U34793 ( .A1(n24903), .A2(n20147), .ZN(n24905) );
OR2_X4 U34794 ( .A1(n20147), .A2(n24903), .ZN(n24904) );
NAND2_X4 U34795 ( .A1(n24905), .A2(n24904), .ZN(n24987) );
NAND2_X4 U34796 ( .A1(n20095), .A2(n24906), .ZN(n24911) );
NAND2_X4 U34797 ( .A1(n20149), .A2(n24907), .ZN(n24909) );
NAND2_X4 U34798 ( .A1(n24909), .A2(n24908), .ZN(n24910) );
NAND2_X4 U34799 ( .A1(n24911), .A2(n24910), .ZN(n24986) );
NOR2_X4 U34800 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_9), .ZN(n24985) );
NOR2_X4 U34801 ( .A1(n24986), .A2(n24985), .ZN(n24912) );
OR2_X4 U34802 ( .A1(n20093), .A2(n24912), .ZN(n24914) );
NAND2_X4 U34803 ( .A1(n24912), .A2(n20093), .ZN(n24913) );
NAND2_X4 U34804 ( .A1(n24914), .A2(n24913), .ZN(n25252) );
NAND2_X4 U34805 ( .A1(n24915), .A2(n24917), .ZN(n24919) );
NAND2_X4 U34806 ( .A1(n24917), .A2(n24916), .ZN(n24918) );
NAND2_X4 U34807 ( .A1(n24919), .A2(n24918), .ZN(n25251) );
NAND2_X4 U34808 ( .A1(n25252), .A2(n25251), .ZN(n24921) );
OR2_X4 U34809 ( .A1(n25251), .A2(n25252), .ZN(n24920) );
NAND2_X4 U34810 ( .A1(n24921), .A2(n24920), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_23_) );
NAND2_X4 U34811 ( .A1(n20148), .A2(n24922), .ZN(n24927) );
NAND2_X4 U34812 ( .A1(n20183), .A2(n24923), .ZN(n24925) );
NAND2_X4 U34813 ( .A1(n24925), .A2(n24924), .ZN(n24926) );
NAND2_X4 U34814 ( .A1(n24927), .A2(n24926), .ZN(n25038) );
NAND2_X4 U34815 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n25037) );
OR2_X4 U34816 ( .A1(n25038), .A2(n20092), .ZN(n24929) );
NAND2_X4 U34817 ( .A1(n20092), .A2(n25038), .ZN(n24928) );
NAND2_X4 U34818 ( .A1(n24929), .A2(n24928), .ZN(n24973) );
NAND2_X4 U34819 ( .A1(n20184), .A2(n20219), .ZN(n24935) );
NAND2_X4 U34820 ( .A1(n24931), .A2(n24930), .ZN(n24933) );
NAND2_X4 U34821 ( .A1(n24933), .A2(n24932), .ZN(n24934) );
NAND2_X4 U34822 ( .A1(n24935), .A2(n24934), .ZN(n24995) );
NAND2_X4 U34823 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n24993) );
OR2_X4 U34824 ( .A1(n24995), .A2(n20146), .ZN(n24937) );
NAND2_X4 U34825 ( .A1(n20146), .A2(n24995), .ZN(n24936) );
NAND2_X4 U34826 ( .A1(n24937), .A2(n24936), .ZN(n24970) );
NAND2_X4 U34827 ( .A1(n20220), .A2(n24938), .ZN(n24943) );
NAND2_X4 U34828 ( .A1(n20255), .A2(n24939), .ZN(n24941) );
NAND2_X4 U34829 ( .A1(n24941), .A2(n24940), .ZN(n24942) );
NAND2_X4 U34830 ( .A1(n24943), .A2(n24942), .ZN(n25003) );
NAND2_X4 U34831 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n25002) );
OR2_X4 U34832 ( .A1(n25003), .A2(n20182), .ZN(n24945) );
NAND2_X4 U34833 ( .A1(n20182), .A2(n25003), .ZN(n24944) );
NAND2_X4 U34834 ( .A1(n24945), .A2(n24944), .ZN(n24967) );
NAND2_X4 U34835 ( .A1(n20256), .A2(n20292), .ZN(n24951) );
NAND2_X4 U34836 ( .A1(n24947), .A2(n24946), .ZN(n24949) );
NAND2_X4 U34837 ( .A1(n24949), .A2(n24948), .ZN(n24950) );
NAND2_X4 U34838 ( .A1(n24951), .A2(n24950), .ZN(n25011) );
NAND2_X4 U34839 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n25009) );
OR2_X4 U34840 ( .A1(n25011), .A2(n20218), .ZN(n24953) );
NAND2_X4 U34841 ( .A1(n20218), .A2(n25011), .ZN(n24952) );
NAND2_X4 U34842 ( .A1(n24953), .A2(n24952), .ZN(n24964) );
NOR2_X4 U34843 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_10), .ZN(n25020) );
NAND2_X4 U34844 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n25019) );
NAND2_X4 U34845 ( .A1(n25020), .A2(n25019), .ZN(n24955) );
OR2_X4 U34846 ( .A1(n25019), .A2(n25020), .ZN(n24954) );
NAND2_X4 U34847 ( .A1(n24955), .A2(n24954), .ZN(n24961) );
NAND2_X4 U34848 ( .A1(n24957), .A2(n20293), .ZN(n24960) );
NAND2_X4 U34849 ( .A1(n20293), .A2(n24958), .ZN(n24959) );
NAND2_X4 U34850 ( .A1(n24960), .A2(n24959), .ZN(n25021) );
NAND2_X4 U34851 ( .A1(n24961), .A2(n25021), .ZN(n24963) );
OR2_X4 U34852 ( .A1(n25021), .A2(n24961), .ZN(n24962) );
NAND2_X4 U34853 ( .A1(n24963), .A2(n24962), .ZN(n25010) );
NAND2_X4 U34854 ( .A1(n24964), .A2(n20253), .ZN(n24966) );
OR2_X4 U34855 ( .A1(n20253), .A2(n24964), .ZN(n24965) );
NAND2_X4 U34856 ( .A1(n24966), .A2(n24965), .ZN(n25001) );
NAND2_X4 U34857 ( .A1(n24967), .A2(n20217), .ZN(n24969) );
OR2_X4 U34858 ( .A1(n20217), .A2(n24967), .ZN(n24968) );
NAND2_X4 U34859 ( .A1(n24969), .A2(n24968), .ZN(n24994) );
NAND2_X4 U34860 ( .A1(n24970), .A2(n20181), .ZN(n24972) );
OR2_X4 U34861 ( .A1(n20181), .A2(n24970), .ZN(n24971) );
NAND2_X4 U34862 ( .A1(n24972), .A2(n24971), .ZN(n25036) );
NAND2_X4 U34863 ( .A1(n24973), .A2(n20145), .ZN(n24975) );
OR2_X4 U34864 ( .A1(n20145), .A2(n24973), .ZN(n24974) );
AND2_X4 U34865 ( .A1(n24975), .A2(n24974), .ZN(n25047) );
NAND2_X4 U34866 ( .A1(n20094), .A2(n20147), .ZN(n24981) );
NAND2_X4 U34867 ( .A1(n24977), .A2(n24976), .ZN(n24979) );
NAND2_X4 U34868 ( .A1(n24979), .A2(n24978), .ZN(n24980) );
NAND2_X4 U34869 ( .A1(n24981), .A2(n24980), .ZN(n25046) );
NOR2_X4 U34870 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_10), .ZN(n25045) );
NOR2_X4 U34871 ( .A1(n25046), .A2(n25045), .ZN(n24982) );
OR2_X4 U34872 ( .A1(n25047), .A2(n24982), .ZN(n24984) );
NAND2_X4 U34873 ( .A1(n24982), .A2(n25047), .ZN(n24983) );
NAND2_X4 U34874 ( .A1(n24984), .A2(n24983), .ZN(n24991) );
NAND2_X4 U34875 ( .A1(n24985), .A2(n24987), .ZN(n24989) );
NAND2_X4 U34876 ( .A1(n24987), .A2(n24986), .ZN(n24988) );
NAND2_X4 U34877 ( .A1(n24989), .A2(n24988), .ZN(n24990) );
NOR2_X4 U34878 ( .A1(n24991), .A2(n24990), .ZN(n24992) );
NOR2_X4 U34879 ( .A1(n20049), .A2(n20048), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_25_) );
NOR2_X4 U34880 ( .A1(n24992), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_25_), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_24_) );
NAND2_X4 U34881 ( .A1(n20146), .A2(n20181), .ZN(n24998) );
NAND2_X4 U34882 ( .A1(n24994), .A2(n24993), .ZN(n24996) );
NAND2_X4 U34883 ( .A1(n24996), .A2(n24995), .ZN(n24997) );
NAND2_X4 U34884 ( .A1(n24998), .A2(n24997), .ZN(n25086) );
NAND2_X4 U34885 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n25084) );
OR2_X4 U34886 ( .A1(n25086), .A2(n20091), .ZN(n25000) );
NAND2_X4 U34887 ( .A1(n20091), .A2(n25086), .ZN(n24999) );
NAND2_X4 U34888 ( .A1(n25000), .A2(n24999), .ZN(n25033) );
NAND2_X4 U34889 ( .A1(n20182), .A2(n25001), .ZN(n25006) );
NAND2_X4 U34890 ( .A1(n20217), .A2(n25002), .ZN(n25004) );
NAND2_X4 U34891 ( .A1(n25004), .A2(n25003), .ZN(n25005) );
NAND2_X4 U34892 ( .A1(n25006), .A2(n25005), .ZN(n25054) );
NAND2_X4 U34893 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n25053) );
OR2_X4 U34894 ( .A1(n25054), .A2(n20144), .ZN(n25008) );
NAND2_X4 U34895 ( .A1(n20144), .A2(n25054), .ZN(n25007) );
NAND2_X4 U34896 ( .A1(n25008), .A2(n25007), .ZN(n25030) );
NAND2_X4 U34897 ( .A1(n20218), .A2(n20253), .ZN(n25014) );
NAND2_X4 U34898 ( .A1(n25010), .A2(n25009), .ZN(n25012) );
NAND2_X4 U34899 ( .A1(n25012), .A2(n25011), .ZN(n25013) );
NAND2_X4 U34900 ( .A1(n25014), .A2(n25013), .ZN(n25062) );
NAND2_X4 U34901 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n25060) );
OR2_X4 U34902 ( .A1(n25062), .A2(n20180), .ZN(n25016) );
NAND2_X4 U34903 ( .A1(n20180), .A2(n25062), .ZN(n25015) );
NAND2_X4 U34904 ( .A1(n25016), .A2(n25015), .ZN(n25027) );
NOR2_X4 U34905 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_11), .ZN(n25071) );
NAND2_X4 U34906 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n25070) );
NAND2_X4 U34907 ( .A1(n25071), .A2(n25070), .ZN(n25018) );
OR2_X4 U34908 ( .A1(n25070), .A2(n25071), .ZN(n25017) );
NAND2_X4 U34909 ( .A1(n25018), .A2(n25017), .ZN(n25024) );
NAND2_X4 U34910 ( .A1(n25020), .A2(n20254), .ZN(n25023) );
NAND2_X4 U34911 ( .A1(n20254), .A2(n25021), .ZN(n25022) );
NAND2_X4 U34912 ( .A1(n25023), .A2(n25022), .ZN(n25072) );
NAND2_X4 U34913 ( .A1(n25024), .A2(n25072), .ZN(n25026) );
OR2_X4 U34914 ( .A1(n25072), .A2(n25024), .ZN(n25025) );
NAND2_X4 U34915 ( .A1(n25026), .A2(n25025), .ZN(n25061) );
NAND2_X4 U34916 ( .A1(n25027), .A2(n20215), .ZN(n25029) );
OR2_X4 U34917 ( .A1(n20215), .A2(n25027), .ZN(n25028) );
NAND2_X4 U34918 ( .A1(n25029), .A2(n25028), .ZN(n25052) );
NAND2_X4 U34919 ( .A1(n25030), .A2(n20179), .ZN(n25032) );
OR2_X4 U34920 ( .A1(n20179), .A2(n25030), .ZN(n25031) );
NAND2_X4 U34921 ( .A1(n25032), .A2(n25031), .ZN(n25085) );
NAND2_X4 U34922 ( .A1(n25033), .A2(n20143), .ZN(n25035) );
OR2_X4 U34923 ( .A1(n20143), .A2(n25033), .ZN(n25034) );
NAND2_X4 U34924 ( .A1(n25035), .A2(n25034), .ZN(n25095) );
NAND2_X4 U34925 ( .A1(n20092), .A2(n25036), .ZN(n25041) );
NAND2_X4 U34926 ( .A1(n20145), .A2(n25037), .ZN(n25039) );
NAND2_X4 U34927 ( .A1(n25039), .A2(n25038), .ZN(n25040) );
NAND2_X4 U34928 ( .A1(n25041), .A2(n25040), .ZN(n25094) );
NOR2_X4 U34929 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_11), .ZN(n25093) );
NOR2_X4 U34930 ( .A1(n25094), .A2(n25093), .ZN(n25042) );
OR2_X4 U34931 ( .A1(n20090), .A2(n25042), .ZN(n25044) );
NAND2_X4 U34932 ( .A1(n25042), .A2(n20090), .ZN(n25043) );
NAND2_X4 U34933 ( .A1(n25044), .A2(n25043), .ZN(n25254) );
NAND2_X4 U34934 ( .A1(n25045), .A2(n25047), .ZN(n25049) );
NAND2_X4 U34935 ( .A1(n25047), .A2(n25046), .ZN(n25048) );
NAND2_X4 U34936 ( .A1(n25049), .A2(n25048), .ZN(n25253) );
NAND2_X4 U34937 ( .A1(n25254), .A2(n25253), .ZN(n25051) );
OR2_X4 U34938 ( .A1(n25253), .A2(n25254), .ZN(n25050) );
NAND2_X4 U34939 ( .A1(n25051), .A2(n25050), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_25_) );
NAND2_X4 U34940 ( .A1(n20144), .A2(n25052), .ZN(n25057) );
NAND2_X4 U34941 ( .A1(n20179), .A2(n25053), .ZN(n25055) );
NAND2_X4 U34942 ( .A1(n25055), .A2(n25054), .ZN(n25056) );
NAND2_X4 U34943 ( .A1(n25057), .A2(n25056), .ZN(n25124) );
NAND2_X4 U34944 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n25123) );
OR2_X4 U34945 ( .A1(n25124), .A2(n20089), .ZN(n25059) );
NAND2_X4 U34946 ( .A1(n20089), .A2(n25124), .ZN(n25058) );
NAND2_X4 U34947 ( .A1(n25059), .A2(n25058), .ZN(n25081) );
NAND2_X4 U34948 ( .A1(n20180), .A2(n20215), .ZN(n25065) );
NAND2_X4 U34949 ( .A1(n25061), .A2(n25060), .ZN(n25063) );
NAND2_X4 U34950 ( .A1(n25063), .A2(n25062), .ZN(n25064) );
NAND2_X4 U34951 ( .A1(n25065), .A2(n25064), .ZN(n25103) );
NAND2_X4 U34952 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n25101) );
OR2_X4 U34953 ( .A1(n25103), .A2(n20142), .ZN(n25067) );
NAND2_X4 U34954 ( .A1(n20142), .A2(n25103), .ZN(n25066) );
NAND2_X4 U34955 ( .A1(n25067), .A2(n25066), .ZN(n25078) );
NOR2_X4 U34956 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_12), .ZN(n25112) );
NAND2_X4 U34957 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n25111) );
NAND2_X4 U34958 ( .A1(n25112), .A2(n25111), .ZN(n25069) );
OR2_X4 U34959 ( .A1(n25111), .A2(n25112), .ZN(n25068) );
NAND2_X4 U34960 ( .A1(n25069), .A2(n25068), .ZN(n25075) );
NAND2_X4 U34961 ( .A1(n25071), .A2(n20216), .ZN(n25074) );
NAND2_X4 U34962 ( .A1(n20216), .A2(n25072), .ZN(n25073) );
NAND2_X4 U34963 ( .A1(n25074), .A2(n25073), .ZN(n25113) );
NAND2_X4 U34964 ( .A1(n25075), .A2(n25113), .ZN(n25077) );
OR2_X4 U34965 ( .A1(n25113), .A2(n25075), .ZN(n25076) );
NAND2_X4 U34966 ( .A1(n25077), .A2(n25076), .ZN(n25102) );
NAND2_X4 U34967 ( .A1(n25078), .A2(n20177), .ZN(n25080) );
OR2_X4 U34968 ( .A1(n20177), .A2(n25078), .ZN(n25079) );
NAND2_X4 U34969 ( .A1(n25080), .A2(n25079), .ZN(n25122) );
NAND2_X4 U34970 ( .A1(n25081), .A2(n20141), .ZN(n25083) );
OR2_X4 U34971 ( .A1(n20141), .A2(n25081), .ZN(n25082) );
AND2_X4 U34972 ( .A1(n25083), .A2(n25082), .ZN(n25133) );
NAND2_X4 U34973 ( .A1(n20091), .A2(n20143), .ZN(n25089) );
NAND2_X4 U34974 ( .A1(n25085), .A2(n25084), .ZN(n25087) );
NAND2_X4 U34975 ( .A1(n25087), .A2(n25086), .ZN(n25088) );
NAND2_X4 U34976 ( .A1(n25089), .A2(n25088), .ZN(n25132) );
NOR2_X4 U34977 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_12), .ZN(n25131) );
NOR2_X4 U34978 ( .A1(n25132), .A2(n25131), .ZN(n25090) );
OR2_X4 U34979 ( .A1(n25133), .A2(n25090), .ZN(n25092) );
NAND2_X4 U34980 ( .A1(n25090), .A2(n25133), .ZN(n25091) );
NAND2_X4 U34981 ( .A1(n25092), .A2(n25091), .ZN(n25099) );
NAND2_X4 U34982 ( .A1(n25093), .A2(n25095), .ZN(n25097) );
NAND2_X4 U34983 ( .A1(n25095), .A2(n25094), .ZN(n25096) );
NAND2_X4 U34984 ( .A1(n25097), .A2(n25096), .ZN(n25098) );
NOR2_X4 U34985 ( .A1(n25099), .A2(n25098), .ZN(n25100) );
NOR2_X4 U34986 ( .A1(n20042), .A2(n20041), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_27_) );
NOR2_X4 U34987 ( .A1(n25100), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_27_), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_26_) );
NAND2_X4 U34988 ( .A1(n20142), .A2(n20177), .ZN(n25106) );
NAND2_X4 U34989 ( .A1(n25102), .A2(n25101), .ZN(n25104) );
NAND2_X4 U34990 ( .A1(n25104), .A2(n25103), .ZN(n25105) );
NAND2_X4 U34991 ( .A1(n25106), .A2(n25105), .ZN(n25150) );
NAND2_X4 U34992 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n25148) );
OR2_X4 U34993 ( .A1(n25150), .A2(n20088), .ZN(n25108) );
NAND2_X4 U34994 ( .A1(n20088), .A2(n25150), .ZN(n25107) );
NAND2_X4 U34995 ( .A1(n25108), .A2(n25107), .ZN(n25119) );
NOR2_X4 U34996 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_13), .ZN(n25141) );
NAND2_X4 U34997 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n25140) );
NAND2_X4 U34998 ( .A1(n25141), .A2(n25140), .ZN(n25110) );
OR2_X4 U34999 ( .A1(n25140), .A2(n25141), .ZN(n25109) );
NAND2_X4 U35000 ( .A1(n25110), .A2(n25109), .ZN(n25116) );
NAND2_X4 U35001 ( .A1(n25112), .A2(n20178), .ZN(n25115) );
NAND2_X4 U35002 ( .A1(n20178), .A2(n25113), .ZN(n25114) );
NAND2_X4 U35003 ( .A1(n25115), .A2(n25114), .ZN(n25142) );
NAND2_X4 U35004 ( .A1(n25116), .A2(n25142), .ZN(n25118) );
OR2_X4 U35005 ( .A1(n25142), .A2(n25116), .ZN(n25117) );
NAND2_X4 U35006 ( .A1(n25118), .A2(n25117), .ZN(n25149) );
NAND2_X4 U35007 ( .A1(n25119), .A2(n20139), .ZN(n25121) );
OR2_X4 U35008 ( .A1(n20139), .A2(n25119), .ZN(n25120) );
NAND2_X4 U35009 ( .A1(n25121), .A2(n25120), .ZN(n25159) );
NAND2_X4 U35010 ( .A1(n20089), .A2(n25122), .ZN(n25127) );
NAND2_X4 U35011 ( .A1(n20141), .A2(n25123), .ZN(n25125) );
NAND2_X4 U35012 ( .A1(n25125), .A2(n25124), .ZN(n25126) );
NAND2_X4 U35013 ( .A1(n25127), .A2(n25126), .ZN(n25158) );
NOR2_X4 U35014 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_13), .ZN(n25157) );
NOR2_X4 U35015 ( .A1(n25158), .A2(n25157), .ZN(n25128) );
OR2_X4 U35016 ( .A1(n20087), .A2(n25128), .ZN(n25130) );
NAND2_X4 U35017 ( .A1(n25128), .A2(n20087), .ZN(n25129) );
NAND2_X4 U35018 ( .A1(n25130), .A2(n25129), .ZN(n25256) );
NAND2_X4 U35019 ( .A1(n25131), .A2(n25133), .ZN(n25135) );
NAND2_X4 U35020 ( .A1(n25133), .A2(n25132), .ZN(n25134) );
NAND2_X4 U35021 ( .A1(n25135), .A2(n25134), .ZN(n25255) );
NAND2_X4 U35022 ( .A1(n25256), .A2(n25255), .ZN(n25137) );
OR2_X4 U35023 ( .A1(n25255), .A2(n25256), .ZN(n25136) );
NAND2_X4 U35024 ( .A1(n25137), .A2(n25136), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_27_) );
NOR2_X4 U35025 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_14), .ZN(n25165) );
NAND2_X4 U35026 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n25166) );
NAND2_X4 U35027 ( .A1(n25165), .A2(n25166), .ZN(n25139) );
OR2_X4 U35028 ( .A1(n25166), .A2(n25165), .ZN(n25138) );
NAND2_X4 U35029 ( .A1(n25139), .A2(n25138), .ZN(n25145) );
NAND2_X4 U35030 ( .A1(n25141), .A2(n20140), .ZN(n25144) );
NAND2_X4 U35031 ( .A1(n20140), .A2(n25142), .ZN(n25143) );
NAND2_X4 U35032 ( .A1(n25144), .A2(n25143), .ZN(n25167) );
NAND2_X4 U35033 ( .A1(n25145), .A2(n25167), .ZN(n25147) );
OR2_X4 U35034 ( .A1(n25145), .A2(n25167), .ZN(n25146) );
AND2_X4 U35035 ( .A1(n25147), .A2(n25146), .ZN(n25177) );
NAND2_X4 U35036 ( .A1(n20088), .A2(n20139), .ZN(n25153) );
NAND2_X4 U35037 ( .A1(n25149), .A2(n25148), .ZN(n25151) );
NAND2_X4 U35038 ( .A1(n25151), .A2(n25150), .ZN(n25152) );
NAND2_X4 U35039 ( .A1(n25153), .A2(n25152), .ZN(n25176) );
NOR2_X4 U35040 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_14), .ZN(n25175) );
NOR2_X4 U35041 ( .A1(n25176), .A2(n25175), .ZN(n25154) );
OR2_X4 U35042 ( .A1(n25177), .A2(n25154), .ZN(n25156) );
NAND2_X4 U35043 ( .A1(n25154), .A2(n25177), .ZN(n25155) );
NAND2_X4 U35044 ( .A1(n25156), .A2(n25155), .ZN(n25163) );
NAND2_X4 U35045 ( .A1(n25157), .A2(n25159), .ZN(n25161) );
NAND2_X4 U35046 ( .A1(n25159), .A2(n25158), .ZN(n25160) );
NAND2_X4 U35047 ( .A1(n25161), .A2(n25160), .ZN(n25162) );
NOR2_X4 U35048 ( .A1(n25163), .A2(n25162), .ZN(n25164) );
NOR2_X4 U35049 ( .A1(n20035), .A2(n20034), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_29_) );
NOR2_X4 U35050 ( .A1(n25164), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_29_), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_28_) );
NOR2_X4 U35051 ( .A1(n25166), .A2(n20138), .ZN(n25168) );
NOR2_X4 U35052 ( .A1(n25168), .A2(n25167), .ZN(n25174) );
NOR2_X4 U35053 ( .A1(n20762), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_15), .ZN(n25169) );
NOR2_X4 U35054 ( .A1(n20084), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_15), .ZN(n25170) );
NOR2_X4 U35055 ( .A1(n25169), .A2(n20030), .ZN(n25172) );
NOR2_X4 U35056 ( .A1(n25170), .A2(n20086), .ZN(n25171) );
NOR2_X4 U35057 ( .A1(n25172), .A2(n25171), .ZN(n25173) );
NAND2_X4 U35058 ( .A1(n25174), .A2(n25173), .ZN(n25181) );
NAND2_X4 U35059 ( .A1(n25175), .A2(n25177), .ZN(n25179) );
NAND2_X4 U35060 ( .A1(n25177), .A2(n25176), .ZN(n25178) );
NAND2_X4 U35061 ( .A1(n25179), .A2(n25178), .ZN(n25180) );
NAND2_X4 U35062 ( .A1(n20029), .A2(n25180), .ZN(n25183) );
NAND2_X4 U35063 ( .A1(n20031), .A2(n25181), .ZN(n25182) );
NAND2_X4 U35064 ( .A1(n25183), .A2(n25182), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_29_) );
NAND2_X4 U35065 ( .A1(n20583), .A2(n25184), .ZN(n25187) );
NAND2_X4 U35066 ( .A1(n20548), .A2(n25185), .ZN(n25186) );
NAND2_X4 U35067 ( .A1(n25187), .A2(n25186), .ZN(n25188) );
NAND2_X4 U35068 ( .A1(n25188), .A2(n20589), .ZN(n25190) );
OR2_X4 U35069 ( .A1(n20589), .A2(n25188), .ZN(n25189) );
NAND2_X4 U35070 ( .A1(n25190), .A2(n25189), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N39) );
NOR2_X4 U35071 ( .A1(n20030), .A2(n20086), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_31_) );
NOR2_X4 U35072 ( .A1(n25192), .A2(n25191), .ZN(n25193) );
NOR2_X4 U35073 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_31_), .A2(n25193), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_30_) );
NAND2_X4 U35074 ( .A1(n20547), .A2(n25194), .ZN(n25197) );
NAND2_X4 U35075 ( .A1(n20510), .A2(n25195), .ZN(n25196) );
NAND2_X4 U35076 ( .A1(n25197), .A2(n25196), .ZN(n25198) );
NOR2_X4 U35077 ( .A1(n25198), .A2(n20551), .ZN(n25200) );
AND2_X4 U35078 ( .A1(n20551), .A2(n25198), .ZN(n25199) );
NOR2_X4 U35079 ( .A1(n25200), .A2(n25199), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N40) );
NAND2_X4 U35080 ( .A1(n20509), .A2(n25201), .ZN(n25204) );
NAND2_X4 U35081 ( .A1(n20472), .A2(n25202), .ZN(n25203) );
NAND2_X4 U35082 ( .A1(n25204), .A2(n25203), .ZN(n25205) );
NAND2_X4 U35083 ( .A1(n25205), .A2(n20513), .ZN(n25207) );
OR2_X4 U35084 ( .A1(n20513), .A2(n25205), .ZN(n25206) );
NAND2_X4 U35085 ( .A1(n25207), .A2(n25206), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N41) );
NAND2_X4 U35086 ( .A1(n20471), .A2(n25208), .ZN(n25211) );
NAND2_X4 U35087 ( .A1(n20434), .A2(n25209), .ZN(n25210) );
NAND2_X4 U35088 ( .A1(n25211), .A2(n25210), .ZN(n25212) );
NOR2_X4 U35089 ( .A1(n25212), .A2(n20475), .ZN(n25214) );
AND2_X4 U35090 ( .A1(n20475), .A2(n25212), .ZN(n25213) );
NOR2_X4 U35091 ( .A1(n25214), .A2(n25213), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N42) );
NAND2_X4 U35092 ( .A1(n20433), .A2(n25215), .ZN(n25218) );
NAND2_X4 U35093 ( .A1(n20397), .A2(n25216), .ZN(n25217) );
NAND2_X4 U35094 ( .A1(n25218), .A2(n25217), .ZN(n25219) );
NAND2_X4 U35095 ( .A1(n25219), .A2(n20437), .ZN(n25221) );
OR2_X4 U35096 ( .A1(n20437), .A2(n25219), .ZN(n25220) );
NAND2_X4 U35097 ( .A1(n25221), .A2(n25220), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N43) );
NAND2_X4 U35098 ( .A1(n20396), .A2(n25222), .ZN(n25225) );
NAND2_X4 U35099 ( .A1(n20360), .A2(n25223), .ZN(n25224) );
NAND2_X4 U35100 ( .A1(n25225), .A2(n25224), .ZN(n25226) );
NOR2_X4 U35101 ( .A1(n25226), .A2(n20400), .ZN(n25228) );
AND2_X4 U35102 ( .A1(n20400), .A2(n25226), .ZN(n25227) );
NOR2_X4 U35103 ( .A1(n25228), .A2(n25227), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N44) );
NAND2_X4 U35104 ( .A1(n20359), .A2(n25229), .ZN(n25232) );
NAND2_X4 U35105 ( .A1(n20323), .A2(n25230), .ZN(n25231) );
NAND2_X4 U35106 ( .A1(n25232), .A2(n25231), .ZN(n25233) );
NAND2_X4 U35107 ( .A1(n25233), .A2(n20363), .ZN(n25235) );
OR2_X4 U35108 ( .A1(n20363), .A2(n25233), .ZN(n25234) );
NAND2_X4 U35109 ( .A1(n25235), .A2(n25234), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N45) );
NAND2_X4 U35110 ( .A1(n20322), .A2(n25236), .ZN(n25239) );
NAND2_X4 U35111 ( .A1(n20286), .A2(n25237), .ZN(n25238) );
NAND2_X4 U35112 ( .A1(n25239), .A2(n25238), .ZN(n25240) );
NOR2_X4 U35113 ( .A1(n25240), .A2(n20324), .ZN(n25242) );
AND2_X4 U35114 ( .A1(n20324), .A2(n25240), .ZN(n25241) );
NOR2_X4 U35115 ( .A1(n25242), .A2(n25241), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N46) );
NAND2_X4 U35116 ( .A1(n25243), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_31_), .ZN(n25244) );
NAND2_X4 U35117 ( .A1(n20081), .A2(n25244), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_15_) );
NOR2_X4 U35118 ( .A1(n20073), .A2(n25246), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_18_) );
NOR2_X4 U35119 ( .A1(n20066), .A2(n25248), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_20_) );
NOR2_X4 U35120 ( .A1(n20059), .A2(n25250), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_22_) );
NOR2_X4 U35121 ( .A1(n20052), .A2(n25252), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_24_) );
NOR2_X4 U35122 ( .A1(n20045), .A2(n25254), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_26_) );
NOR2_X4 U35123 ( .A1(n20038), .A2(n25256), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_28_) );
NOR2_X4 U35124 ( .A1(n20031), .A2(n20029), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_30_) );
NOR2_X4 U35125 ( .A1(n20807), .A2(n16200), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N35) );
NAND2_X4 U35126 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_b_1), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_gen_mult_fast_mult_op_a_0), .ZN(n25257) );
OR2_X4 U35127 ( .A1(n25257), .A2(n25258), .ZN(n25260) );
NAND2_X4 U35128 ( .A1(n25258), .A2(n25257), .ZN(n25259) );
NAND2_X4 U35129 ( .A1(n25260), .A2(n25259), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N36) );
NOR2_X4 U35130 ( .A1(n25261), .A2(n25262), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N68) );
AND2_X4 U35131 ( .A1(n25263), .A2(n25264), .ZN(n25262) );
NOR2_X4 U35132 ( .A1(n25264), .A2(n25263), .ZN(n25261) );
NAND2_X4 U35133 ( .A1(n25265), .A2(n25266), .ZN(n25263) );
NAND2_X4 U35134 ( .A1(n25267), .A2(n25268), .ZN(n25266) );
NAND2_X4 U35135 ( .A1(n25269), .A2(n25270), .ZN(n25264) );
NAND2_X4 U35136 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_31_), .A2(n20080), .ZN(n25270) );
OR2_X4 U35137 ( .A1(n20080), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_31_), .ZN(n25269) );
NOR2_X4 U35138 ( .A1(n25271), .A2(n25272), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N67) );
NOR2_X4 U35139 ( .A1(n20028), .A2(n25273), .ZN(n25272) );
AND2_X4 U35140 ( .A1(n25273), .A2(n20028), .ZN(n25271) );
NAND2_X4 U35141 ( .A1(n25274), .A2(n25275), .ZN(n25267) );
NAND2_X4 U35142 ( .A1(n25276), .A2(n25277), .ZN(n25275) );
NAND2_X4 U35143 ( .A1(n25268), .A2(n25265), .ZN(n25273) );
NAND2_X4 U35144 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_30_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_30_), .ZN(n25265) );
OR2_X4 U35145 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_30_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_30_), .ZN(n25268) );
NOR2_X4 U35146 ( .A1(n25278), .A2(n25279), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N66) );
NOR2_X4 U35147 ( .A1(n20033), .A2(n25280), .ZN(n25279) );
AND2_X4 U35148 ( .A1(n25280), .A2(n20033), .ZN(n25278) );
NAND2_X4 U35149 ( .A1(n25281), .A2(n25282), .ZN(n25276) );
NAND2_X4 U35150 ( .A1(n25283), .A2(n25284), .ZN(n25282) );
NAND2_X4 U35151 ( .A1(n25277), .A2(n25274), .ZN(n25280) );
NAND2_X4 U35152 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_29_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_29_), .ZN(n25274) );
OR2_X4 U35153 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_29_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_29_), .ZN(n25277) );
NOR2_X4 U35154 ( .A1(n25285), .A2(n25286), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N65) );
NOR2_X4 U35155 ( .A1(n20037), .A2(n25287), .ZN(n25286) );
AND2_X4 U35156 ( .A1(n25287), .A2(n20037), .ZN(n25285) );
NAND2_X4 U35157 ( .A1(n25288), .A2(n25289), .ZN(n25283) );
NAND2_X4 U35158 ( .A1(n25290), .A2(n25291), .ZN(n25289) );
NAND2_X4 U35159 ( .A1(n25284), .A2(n25281), .ZN(n25287) );
NAND2_X4 U35160 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_28_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_28_), .ZN(n25281) );
OR2_X4 U35161 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_28_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_28_), .ZN(n25284) );
NOR2_X4 U35162 ( .A1(n25292), .A2(n25293), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N64) );
NOR2_X4 U35163 ( .A1(n20040), .A2(n25294), .ZN(n25293) );
AND2_X4 U35164 ( .A1(n25294), .A2(n20040), .ZN(n25292) );
NAND2_X4 U35165 ( .A1(n25295), .A2(n25296), .ZN(n25290) );
NAND2_X4 U35166 ( .A1(n25297), .A2(n25298), .ZN(n25296) );
NAND2_X4 U35167 ( .A1(n25291), .A2(n25288), .ZN(n25294) );
NAND2_X4 U35168 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_27_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_27_), .ZN(n25288) );
OR2_X4 U35169 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_27_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_27_), .ZN(n25291) );
NOR2_X4 U35170 ( .A1(n25299), .A2(n25300), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N63) );
NOR2_X4 U35171 ( .A1(n20044), .A2(n25301), .ZN(n25300) );
AND2_X4 U35172 ( .A1(n25301), .A2(n20044), .ZN(n25299) );
NAND2_X4 U35173 ( .A1(n25302), .A2(n25303), .ZN(n25297) );
NAND2_X4 U35174 ( .A1(n25304), .A2(n25305), .ZN(n25303) );
NAND2_X4 U35175 ( .A1(n25298), .A2(n25295), .ZN(n25301) );
NAND2_X4 U35176 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_26_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_26_), .ZN(n25295) );
OR2_X4 U35177 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_26_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_26_), .ZN(n25298) );
NOR2_X4 U35178 ( .A1(n25306), .A2(n25307), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N62) );
NOR2_X4 U35179 ( .A1(n20047), .A2(n25308), .ZN(n25307) );
AND2_X4 U35180 ( .A1(n25308), .A2(n20047), .ZN(n25306) );
NAND2_X4 U35181 ( .A1(n25309), .A2(n25310), .ZN(n25304) );
NAND2_X4 U35182 ( .A1(n25311), .A2(n25312), .ZN(n25310) );
NAND2_X4 U35183 ( .A1(n25305), .A2(n25302), .ZN(n25308) );
NAND2_X4 U35184 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_25_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_25_), .ZN(n25302) );
OR2_X4 U35185 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_25_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_25_), .ZN(n25305) );
NOR2_X4 U35186 ( .A1(n25313), .A2(n25314), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N61) );
NOR2_X4 U35187 ( .A1(n20051), .A2(n25315), .ZN(n25314) );
AND2_X4 U35188 ( .A1(n25315), .A2(n20051), .ZN(n25313) );
NAND2_X4 U35189 ( .A1(n25316), .A2(n25317), .ZN(n25311) );
NAND2_X4 U35190 ( .A1(n25318), .A2(n25319), .ZN(n25317) );
NAND2_X4 U35191 ( .A1(n25312), .A2(n25309), .ZN(n25315) );
NAND2_X4 U35192 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_24_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_24_), .ZN(n25309) );
OR2_X4 U35193 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_24_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_24_), .ZN(n25312) );
NOR2_X4 U35194 ( .A1(n25320), .A2(n25321), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N60) );
NOR2_X4 U35195 ( .A1(n20054), .A2(n25322), .ZN(n25321) );
AND2_X4 U35196 ( .A1(n25322), .A2(n20054), .ZN(n25320) );
NAND2_X4 U35197 ( .A1(n25323), .A2(n25324), .ZN(n25318) );
NAND2_X4 U35198 ( .A1(n25325), .A2(n25326), .ZN(n25324) );
NAND2_X4 U35199 ( .A1(n25319), .A2(n25316), .ZN(n25322) );
NAND2_X4 U35200 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_23_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_23_), .ZN(n25316) );
OR2_X4 U35201 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_23_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_23_), .ZN(n25319) );
NOR2_X4 U35202 ( .A1(n25327), .A2(n25328), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N59) );
NOR2_X4 U35203 ( .A1(n20058), .A2(n25329), .ZN(n25328) );
AND2_X4 U35204 ( .A1(n25329), .A2(n20058), .ZN(n25327) );
NAND2_X4 U35205 ( .A1(n25330), .A2(n25331), .ZN(n25325) );
NAND2_X4 U35206 ( .A1(n25332), .A2(n25333), .ZN(n25331) );
NAND2_X4 U35207 ( .A1(n25326), .A2(n25323), .ZN(n25329) );
NAND2_X4 U35208 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_22_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_22_), .ZN(n25323) );
OR2_X4 U35209 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_22_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_22_), .ZN(n25326) );
NOR2_X4 U35210 ( .A1(n25334), .A2(n25335), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N58) );
NOR2_X4 U35211 ( .A1(n20061), .A2(n25336), .ZN(n25335) );
AND2_X4 U35212 ( .A1(n25336), .A2(n20061), .ZN(n25334) );
NAND2_X4 U35213 ( .A1(n25337), .A2(n25338), .ZN(n25332) );
NAND2_X4 U35214 ( .A1(n25339), .A2(n25340), .ZN(n25338) );
NAND2_X4 U35215 ( .A1(n25333), .A2(n25330), .ZN(n25336) );
NAND2_X4 U35216 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_21_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_21_), .ZN(n25330) );
OR2_X4 U35217 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_21_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_21_), .ZN(n25333) );
NOR2_X4 U35218 ( .A1(n25341), .A2(n25342), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N57) );
NOR2_X4 U35219 ( .A1(n20065), .A2(n25343), .ZN(n25342) );
AND2_X4 U35220 ( .A1(n25343), .A2(n20065), .ZN(n25341) );
NAND2_X4 U35221 ( .A1(n25344), .A2(n25345), .ZN(n25339) );
NAND2_X4 U35222 ( .A1(n25346), .A2(n25347), .ZN(n25345) );
NAND2_X4 U35223 ( .A1(n25340), .A2(n25337), .ZN(n25343) );
NAND2_X4 U35224 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_20_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_20_), .ZN(n25337) );
OR2_X4 U35225 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_20_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_20_), .ZN(n25340) );
NOR2_X4 U35226 ( .A1(n25348), .A2(n25349), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N56) );
NOR2_X4 U35227 ( .A1(n20068), .A2(n25350), .ZN(n25349) );
AND2_X4 U35228 ( .A1(n25350), .A2(n20068), .ZN(n25348) );
NAND2_X4 U35229 ( .A1(n25351), .A2(n25352), .ZN(n25346) );
NAND2_X4 U35230 ( .A1(n25353), .A2(n25354), .ZN(n25352) );
NAND2_X4 U35231 ( .A1(n25347), .A2(n25344), .ZN(n25350) );
NAND2_X4 U35232 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_19_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_19_), .ZN(n25344) );
OR2_X4 U35233 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_19_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_19_), .ZN(n25347) );
NOR2_X4 U35234 ( .A1(n25355), .A2(n25356), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N55) );
NOR2_X4 U35235 ( .A1(n20072), .A2(n25357), .ZN(n25356) );
AND2_X4 U35236 ( .A1(n25357), .A2(n20072), .ZN(n25355) );
NAND2_X4 U35237 ( .A1(n25358), .A2(n25359), .ZN(n25353) );
NAND2_X4 U35238 ( .A1(n25360), .A2(n25361), .ZN(n25359) );
NAND2_X4 U35239 ( .A1(n25354), .A2(n25351), .ZN(n25357) );
NAND2_X4 U35240 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_18_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_18_), .ZN(n25351) );
OR2_X4 U35241 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_18_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_18_), .ZN(n25354) );
NOR2_X4 U35242 ( .A1(n25362), .A2(n25363), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N54) );
NOR2_X4 U35243 ( .A1(n20075), .A2(n25364), .ZN(n25363) );
AND2_X4 U35244 ( .A1(n25364), .A2(n20075), .ZN(n25362) );
NAND2_X4 U35245 ( .A1(n25365), .A2(n25366), .ZN(n25360) );
NAND2_X4 U35246 ( .A1(n25367), .A2(n25368), .ZN(n25366) );
NAND2_X4 U35247 ( .A1(n25361), .A2(n25358), .ZN(n25364) );
NAND2_X4 U35248 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_17_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_17_), .ZN(n25358) );
OR2_X4 U35249 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_17_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_17_), .ZN(n25361) );
NAND2_X4 U35250 ( .A1(n25369), .A2(n25370), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N53) );
NAND2_X4 U35251 ( .A1(n25367), .A2(n25371), .ZN(n25370) );
OR2_X4 U35252 ( .A1(n25371), .A2(n25367), .ZN(n25369) );
NAND2_X4 U35253 ( .A1(n25368), .A2(n25365), .ZN(n25371) );
NAND2_X4 U35254 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_16_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_16_), .ZN(n25365) );
OR2_X4 U35255 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_16_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_16_), .ZN(n25368) );
NOR2_X4 U35256 ( .A1(n25367), .A2(n25372), .ZN(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N52) );
NOR2_X4 U35257 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_15_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_15_), .ZN(n25372) );
AND2_X4 U35258 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A2_15_), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_mult_268_A1_15_), .ZN(n25367) );
OR2_X4 U35259 ( .A1(n20682), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_0), .ZN(n25374) );
NAND2_X4 U35260 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_0), .A2(n20682), .ZN(n25373) );
NAND2_X4 U35261 ( .A1(n25374), .A2(n25373), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_0) );
NAND2_X4 U35262 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_0), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N35), .ZN(n25490) );
OR2_X4 U35263 ( .A1(n20673), .A2(n25490), .ZN(n25377) );
NAND2_X4 U35264 ( .A1(n20673), .A2(n25490), .ZN(n25375) );
NAND2_X4 U35265 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_1), .A2(n25375), .ZN(n25376) );
NAND2_X4 U35266 ( .A1(n25377), .A2(n25376), .ZN(n25587) );
NAND2_X4 U35267 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N37), .A2(n25587), .ZN(n25380) );
OR2_X4 U35268 ( .A1(n25587), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N37), .ZN(n25378) );
NAND2_X4 U35269 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_2), .A2(n25378), .ZN(n25379) );
NAND2_X4 U35270 ( .A1(n25380), .A2(n25379), .ZN(n25630) );
NAND2_X4 U35271 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N38), .A2(n25630), .ZN(n25383) );
OR2_X4 U35272 ( .A1(n25630), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N38), .ZN(n25381) );
NAND2_X4 U35273 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_3), .A2(n25381), .ZN(n25382) );
NAND2_X4 U35274 ( .A1(n25383), .A2(n25382), .ZN(n25636) );
NAND2_X4 U35275 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N39), .A2(n25636), .ZN(n25386) );
OR2_X4 U35276 ( .A1(n25636), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N39), .ZN(n25384) );
NAND2_X4 U35277 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_4), .A2(n25384), .ZN(n25385) );
NAND2_X4 U35278 ( .A1(n25386), .A2(n25385), .ZN(n25642) );
NAND2_X4 U35279 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N40), .A2(n25642), .ZN(n25389) );
OR2_X4 U35280 ( .A1(n25642), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N40), .ZN(n25387) );
NAND2_X4 U35281 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_5), .A2(n25387), .ZN(n25388) );
NAND2_X4 U35282 ( .A1(n25389), .A2(n25388), .ZN(n25648) );
NAND2_X4 U35283 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N41), .A2(n25648), .ZN(n25392) );
OR2_X4 U35284 ( .A1(n25648), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N41), .ZN(n25390) );
NAND2_X4 U35285 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_6), .A2(n25390), .ZN(n25391) );
NAND2_X4 U35286 ( .A1(n25392), .A2(n25391), .ZN(n25654) );
NAND2_X4 U35287 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N42), .A2(n25654), .ZN(n25395) );
OR2_X4 U35288 ( .A1(n25654), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N42), .ZN(n25393) );
NAND2_X4 U35289 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_7), .A2(n25393), .ZN(n25394) );
NAND2_X4 U35290 ( .A1(n25395), .A2(n25394), .ZN(n25660) );
NAND2_X4 U35291 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N43), .A2(n25660), .ZN(n25398) );
OR2_X4 U35292 ( .A1(n25660), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N43), .ZN(n25396) );
NAND2_X4 U35293 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_8), .A2(n25396), .ZN(n25397) );
NAND2_X4 U35294 ( .A1(n25398), .A2(n25397), .ZN(n25666) );
NAND2_X4 U35295 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N44), .A2(n25666), .ZN(n25401) );
OR2_X4 U35296 ( .A1(n25666), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N44), .ZN(n25399) );
NAND2_X4 U35297 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_9), .A2(n25399), .ZN(n25400) );
NAND2_X4 U35298 ( .A1(n25401), .A2(n25400), .ZN(n25407) );
OR2_X4 U35299 ( .A1(n20321), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_10), .ZN(n25403) );
NAND2_X4 U35300 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_10), .A2(n20321), .ZN(n25402) );
NAND2_X4 U35301 ( .A1(n25403), .A2(n25402), .ZN(n25404) );
NOR2_X4 U35302 ( .A1(n25407), .A2(n25404), .ZN(n25406) );
AND2_X4 U35303 ( .A1(n25407), .A2(n25404), .ZN(n25405) );
NOR2_X4 U35304 ( .A1(n25406), .A2(n25405), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_10) );
NAND2_X4 U35305 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N45), .A2(n25407), .ZN(n25410) );
OR2_X4 U35306 ( .A1(n25407), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N45), .ZN(n25408) );
NAND2_X4 U35307 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_10), .A2(n25408), .ZN(n25409) );
NAND2_X4 U35308 ( .A1(n25410), .A2(n25409), .ZN(n25416) );
OR2_X4 U35309 ( .A1(n20284), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_11), .ZN(n25412) );
NAND2_X4 U35310 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_11), .A2(n20284), .ZN(n25411) );
NAND2_X4 U35311 ( .A1(n25412), .A2(n25411), .ZN(n25413) );
NOR2_X4 U35312 ( .A1(n25416), .A2(n25413), .ZN(n25415) );
AND2_X4 U35313 ( .A1(n25416), .A2(n25413), .ZN(n25414) );
NOR2_X4 U35314 ( .A1(n25415), .A2(n25414), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_11) );
NAND2_X4 U35315 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N46), .A2(n25416), .ZN(n25419) );
OR2_X4 U35316 ( .A1(n25416), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N46), .ZN(n25417) );
NAND2_X4 U35317 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_11), .A2(n25417), .ZN(n25418) );
NAND2_X4 U35318 ( .A1(n25419), .A2(n25418), .ZN(n25425) );
OR2_X4 U35319 ( .A1(n20246), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_12), .ZN(n25421) );
NAND2_X4 U35320 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_12), .A2(n20246), .ZN(n25420) );
NAND2_X4 U35321 ( .A1(n25421), .A2(n25420), .ZN(n25422) );
NOR2_X4 U35322 ( .A1(n25425), .A2(n25422), .ZN(n25424) );
AND2_X4 U35323 ( .A1(n25425), .A2(n25422), .ZN(n25423) );
NOR2_X4 U35324 ( .A1(n25424), .A2(n25423), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_12) );
NAND2_X4 U35325 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N47), .A2(n25425), .ZN(n25428) );
OR2_X4 U35326 ( .A1(n25425), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N47), .ZN(n25426) );
NAND2_X4 U35327 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_12), .A2(n25426), .ZN(n25427) );
NAND2_X4 U35328 ( .A1(n25428), .A2(n25427), .ZN(n25434) );
OR2_X4 U35329 ( .A1(n20208), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_13), .ZN(n25430) );
NAND2_X4 U35330 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_13), .A2(n20208), .ZN(n25429) );
NAND2_X4 U35331 ( .A1(n25430), .A2(n25429), .ZN(n25431) );
NOR2_X4 U35332 ( .A1(n25434), .A2(n25431), .ZN(n25433) );
AND2_X4 U35333 ( .A1(n25434), .A2(n25431), .ZN(n25432) );
NOR2_X4 U35334 ( .A1(n25433), .A2(n25432), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_13) );
NAND2_X4 U35335 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N48), .A2(n25434), .ZN(n25437) );
OR2_X4 U35336 ( .A1(n25434), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N48), .ZN(n25435) );
NAND2_X4 U35337 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_13), .A2(n25435), .ZN(n25436) );
NAND2_X4 U35338 ( .A1(n25437), .A2(n25436), .ZN(n25443) );
OR2_X4 U35339 ( .A1(n20170), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_14), .ZN(n25439) );
NAND2_X4 U35340 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_14), .A2(n20170), .ZN(n25438) );
NAND2_X4 U35341 ( .A1(n25439), .A2(n25438), .ZN(n25440) );
NOR2_X4 U35342 ( .A1(n25443), .A2(n25440), .ZN(n25442) );
AND2_X4 U35343 ( .A1(n25443), .A2(n25440), .ZN(n25441) );
NOR2_X4 U35344 ( .A1(n25442), .A2(n25441), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_14) );
NAND2_X4 U35345 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N49), .A2(n25443), .ZN(n25446) );
OR2_X4 U35346 ( .A1(n25443), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N49), .ZN(n25444) );
NAND2_X4 U35347 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_14), .A2(n25444), .ZN(n25445) );
NAND2_X4 U35348 ( .A1(n25446), .A2(n25445), .ZN(n25452) );
OR2_X4 U35349 ( .A1(n20108), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_15), .ZN(n25448) );
NAND2_X4 U35350 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_15), .A2(n20108), .ZN(n25447) );
NAND2_X4 U35351 ( .A1(n25448), .A2(n25447), .ZN(n25449) );
NOR2_X4 U35352 ( .A1(n25452), .A2(n25449), .ZN(n25451) );
AND2_X4 U35353 ( .A1(n25452), .A2(n25449), .ZN(n25450) );
NOR2_X4 U35354 ( .A1(n25451), .A2(n25450), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_15) );
NAND2_X4 U35355 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N50), .A2(n25452), .ZN(n25455) );
OR2_X4 U35356 ( .A1(n25452), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N50), .ZN(n25453) );
NAND2_X4 U35357 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_15), .A2(n25453), .ZN(n25454) );
NAND2_X4 U35358 ( .A1(n25455), .A2(n25454), .ZN(n25461) );
OR2_X4 U35359 ( .A1(n20026), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_16), .ZN(n25457) );
NAND2_X4 U35360 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_16), .A2(n20026), .ZN(n25456) );
NAND2_X4 U35361 ( .A1(n25457), .A2(n25456), .ZN(n25458) );
NOR2_X4 U35362 ( .A1(n25461), .A2(n25458), .ZN(n25460) );
AND2_X4 U35363 ( .A1(n25461), .A2(n25458), .ZN(n25459) );
NOR2_X4 U35364 ( .A1(n25460), .A2(n25459), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_16) );
NAND2_X4 U35365 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N51), .A2(n25461), .ZN(n25464) );
OR2_X4 U35366 ( .A1(n25461), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N51), .ZN(n25462) );
NAND2_X4 U35367 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_16), .A2(n25462), .ZN(n25463) );
NAND2_X4 U35368 ( .A1(n25464), .A2(n25463), .ZN(n25470) );
OR2_X4 U35369 ( .A1(n20078), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_17), .ZN(n25466) );
NAND2_X4 U35370 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_17), .A2(n20078), .ZN(n25465) );
NAND2_X4 U35371 ( .A1(n25466), .A2(n25465), .ZN(n25467) );
NOR2_X4 U35372 ( .A1(n25470), .A2(n25467), .ZN(n25469) );
AND2_X4 U35373 ( .A1(n25470), .A2(n25467), .ZN(n25468) );
NOR2_X4 U35374 ( .A1(n25469), .A2(n25468), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_17) );
NAND2_X4 U35375 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N52), .A2(n25470), .ZN(n25473) );
OR2_X4 U35376 ( .A1(n25470), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N52), .ZN(n25471) );
NAND2_X4 U35377 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_17), .A2(n25471), .ZN(n25472) );
NAND2_X4 U35378 ( .A1(n25473), .A2(n25472), .ZN(n25479) );
OR2_X4 U35379 ( .A1(n20074), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_18), .ZN(n25475) );
NAND2_X4 U35380 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_18), .A2(n20074), .ZN(n25474) );
NAND2_X4 U35381 ( .A1(n25475), .A2(n25474), .ZN(n25476) );
NOR2_X4 U35382 ( .A1(n25479), .A2(n25476), .ZN(n25478) );
AND2_X4 U35383 ( .A1(n25479), .A2(n25476), .ZN(n25477) );
NOR2_X4 U35384 ( .A1(n25478), .A2(n25477), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_18) );
NAND2_X4 U35385 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N53), .A2(n25479), .ZN(n25482) );
OR2_X4 U35386 ( .A1(n25479), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N53), .ZN(n25480) );
NAND2_X4 U35387 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_18), .A2(n25480), .ZN(n25481) );
NAND2_X4 U35388 ( .A1(n25482), .A2(n25481), .ZN(n25494) );
OR2_X4 U35389 ( .A1(n20071), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_19), .ZN(n25484) );
NAND2_X4 U35390 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_19), .A2(n20071), .ZN(n25483) );
NAND2_X4 U35391 ( .A1(n25484), .A2(n25483), .ZN(n25485) );
NOR2_X4 U35392 ( .A1(n25494), .A2(n25485), .ZN(n25487) );
AND2_X4 U35393 ( .A1(n25494), .A2(n25485), .ZN(n25486) );
NOR2_X4 U35394 ( .A1(n25487), .A2(n25486), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_19) );
OR2_X4 U35395 ( .A1(n20673), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_1), .ZN(n25489) );
NAND2_X4 U35396 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_1), .A2(n20673), .ZN(n25488) );
NAND2_X4 U35397 ( .A1(n25489), .A2(n25488), .ZN(n25491) );
NAND2_X4 U35398 ( .A1(n25491), .A2(n25490), .ZN(n25493) );
OR2_X4 U35399 ( .A1(n25491), .A2(n25490), .ZN(n25492) );
NAND2_X4 U35400 ( .A1(n25493), .A2(n25492), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_1) );
NAND2_X4 U35401 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N54), .A2(n25494), .ZN(n25497) );
OR2_X4 U35402 ( .A1(n25494), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N54), .ZN(n25495) );
NAND2_X4 U35403 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_19), .A2(n25495), .ZN(n25496) );
NAND2_X4 U35404 ( .A1(n25497), .A2(n25496), .ZN(n25503) );
OR2_X4 U35405 ( .A1(n20067), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_20), .ZN(n25499) );
NAND2_X4 U35406 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_20), .A2(n20067), .ZN(n25498) );
NAND2_X4 U35407 ( .A1(n25499), .A2(n25498), .ZN(n25500) );
NOR2_X4 U35408 ( .A1(n25503), .A2(n25500), .ZN(n25502) );
AND2_X4 U35409 ( .A1(n25503), .A2(n25500), .ZN(n25501) );
NOR2_X4 U35410 ( .A1(n25502), .A2(n25501), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_20) );
NAND2_X4 U35411 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N55), .A2(n25503), .ZN(n25506) );
OR2_X4 U35412 ( .A1(n25503), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N55), .ZN(n25504) );
NAND2_X4 U35413 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_20), .A2(n25504), .ZN(n25505) );
NAND2_X4 U35414 ( .A1(n25506), .A2(n25505), .ZN(n25512) );
OR2_X4 U35415 ( .A1(n20064), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_21), .ZN(n25508) );
NAND2_X4 U35416 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_21), .A2(n20064), .ZN(n25507) );
NAND2_X4 U35417 ( .A1(n25508), .A2(n25507), .ZN(n25509) );
NOR2_X4 U35418 ( .A1(n25512), .A2(n25509), .ZN(n25511) );
AND2_X4 U35419 ( .A1(n25512), .A2(n25509), .ZN(n25510) );
NOR2_X4 U35420 ( .A1(n25511), .A2(n25510), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_21) );
NAND2_X4 U35421 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N56), .A2(n25512), .ZN(n25515) );
OR2_X4 U35422 ( .A1(n25512), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N56), .ZN(n25513) );
NAND2_X4 U35423 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_21), .A2(n25513), .ZN(n25514) );
NAND2_X4 U35424 ( .A1(n25515), .A2(n25514), .ZN(n25521) );
OR2_X4 U35425 ( .A1(n20060), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_22), .ZN(n25517) );
NAND2_X4 U35426 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_22), .A2(n20060), .ZN(n25516) );
NAND2_X4 U35427 ( .A1(n25517), .A2(n25516), .ZN(n25518) );
NOR2_X4 U35428 ( .A1(n25521), .A2(n25518), .ZN(n25520) );
AND2_X4 U35429 ( .A1(n25521), .A2(n25518), .ZN(n25519) );
NOR2_X4 U35430 ( .A1(n25520), .A2(n25519), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_22) );
NAND2_X4 U35431 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N57), .A2(n25521), .ZN(n25524) );
OR2_X4 U35432 ( .A1(n25521), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N57), .ZN(n25522) );
NAND2_X4 U35433 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_22), .A2(n25522), .ZN(n25523) );
NAND2_X4 U35434 ( .A1(n25524), .A2(n25523), .ZN(n25530) );
OR2_X4 U35435 ( .A1(n20057), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_23), .ZN(n25526) );
NAND2_X4 U35436 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_23), .A2(n20057), .ZN(n25525) );
NAND2_X4 U35437 ( .A1(n25526), .A2(n25525), .ZN(n25527) );
NOR2_X4 U35438 ( .A1(n25530), .A2(n25527), .ZN(n25529) );
AND2_X4 U35439 ( .A1(n25530), .A2(n25527), .ZN(n25528) );
NOR2_X4 U35440 ( .A1(n25529), .A2(n25528), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_23) );
NAND2_X4 U35441 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N58), .A2(n25530), .ZN(n25533) );
OR2_X4 U35442 ( .A1(n25530), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N58), .ZN(n25531) );
NAND2_X4 U35443 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_23), .A2(n25531), .ZN(n25532) );
NAND2_X4 U35444 ( .A1(n25533), .A2(n25532), .ZN(n25539) );
OR2_X4 U35445 ( .A1(n20053), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_24), .ZN(n25535) );
NAND2_X4 U35446 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_24), .A2(n20053), .ZN(n25534) );
NAND2_X4 U35447 ( .A1(n25535), .A2(n25534), .ZN(n25536) );
NOR2_X4 U35448 ( .A1(n25539), .A2(n25536), .ZN(n25538) );
AND2_X4 U35449 ( .A1(n25539), .A2(n25536), .ZN(n25537) );
NOR2_X4 U35450 ( .A1(n25538), .A2(n25537), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_24) );
NAND2_X4 U35451 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N59), .A2(n25539), .ZN(n25542) );
OR2_X4 U35452 ( .A1(n25539), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N59), .ZN(n25540) );
NAND2_X4 U35453 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_24), .A2(n25540), .ZN(n25541) );
NAND2_X4 U35454 ( .A1(n25542), .A2(n25541), .ZN(n25548) );
OR2_X4 U35455 ( .A1(n20050), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_25), .ZN(n25544) );
NAND2_X4 U35456 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_25), .A2(n20050), .ZN(n25543) );
NAND2_X4 U35457 ( .A1(n25544), .A2(n25543), .ZN(n25545) );
NOR2_X4 U35458 ( .A1(n25548), .A2(n25545), .ZN(n25547) );
AND2_X4 U35459 ( .A1(n25548), .A2(n25545), .ZN(n25546) );
NOR2_X4 U35460 ( .A1(n25547), .A2(n25546), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_25) );
NAND2_X4 U35461 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N60), .A2(n25548), .ZN(n25551) );
OR2_X4 U35462 ( .A1(n25548), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N60), .ZN(n25549) );
NAND2_X4 U35463 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_25), .A2(n25549), .ZN(n25550) );
NAND2_X4 U35464 ( .A1(n25551), .A2(n25550), .ZN(n25557) );
OR2_X4 U35465 ( .A1(n20046), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_26), .ZN(n25553) );
NAND2_X4 U35466 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_26), .A2(n20046), .ZN(n25552) );
NAND2_X4 U35467 ( .A1(n25553), .A2(n25552), .ZN(n25554) );
NOR2_X4 U35468 ( .A1(n25557), .A2(n25554), .ZN(n25556) );
AND2_X4 U35469 ( .A1(n25557), .A2(n25554), .ZN(n25555) );
NOR2_X4 U35470 ( .A1(n25556), .A2(n25555), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_26) );
NAND2_X4 U35471 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N61), .A2(n25557), .ZN(n25560) );
OR2_X4 U35472 ( .A1(n25557), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N61), .ZN(n25558) );
NAND2_X4 U35473 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_26), .A2(n25558), .ZN(n25559) );
NAND2_X4 U35474 ( .A1(n25560), .A2(n25559), .ZN(n25566) );
OR2_X4 U35475 ( .A1(n20043), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_27), .ZN(n25562) );
NAND2_X4 U35476 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_27), .A2(n20043), .ZN(n25561) );
NAND2_X4 U35477 ( .A1(n25562), .A2(n25561), .ZN(n25563) );
NOR2_X4 U35478 ( .A1(n25566), .A2(n25563), .ZN(n25565) );
AND2_X4 U35479 ( .A1(n25566), .A2(n25563), .ZN(n25564) );
NOR2_X4 U35480 ( .A1(n25565), .A2(n25564), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_27) );
NAND2_X4 U35481 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N62), .A2(n25566), .ZN(n25569) );
OR2_X4 U35482 ( .A1(n25566), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N62), .ZN(n25567) );
NAND2_X4 U35483 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_27), .A2(n25567), .ZN(n25568) );
NAND2_X4 U35484 ( .A1(n25569), .A2(n25568), .ZN(n25575) );
OR2_X4 U35485 ( .A1(n20039), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_28), .ZN(n25571) );
NAND2_X4 U35486 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_28), .A2(n20039), .ZN(n25570) );
NAND2_X4 U35487 ( .A1(n25571), .A2(n25570), .ZN(n25572) );
NOR2_X4 U35488 ( .A1(n25575), .A2(n25572), .ZN(n25574) );
AND2_X4 U35489 ( .A1(n25575), .A2(n25572), .ZN(n25573) );
NOR2_X4 U35490 ( .A1(n25574), .A2(n25573), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_28) );
NAND2_X4 U35491 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N63), .A2(n25575), .ZN(n25578) );
OR2_X4 U35492 ( .A1(n25575), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N63), .ZN(n25576) );
NAND2_X4 U35493 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_28), .A2(n25576), .ZN(n25577) );
NAND2_X4 U35494 ( .A1(n25578), .A2(n25577), .ZN(n25590) );
OR2_X4 U35495 ( .A1(n20036), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_29), .ZN(n25580) );
NAND2_X4 U35496 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_29), .A2(n20036), .ZN(n25579) );
NAND2_X4 U35497 ( .A1(n25580), .A2(n25579), .ZN(n25581) );
NOR2_X4 U35498 ( .A1(n25590), .A2(n25581), .ZN(n25583) );
AND2_X4 U35499 ( .A1(n25590), .A2(n25581), .ZN(n25582) );
NOR2_X4 U35500 ( .A1(n25583), .A2(n25582), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_29) );
OR2_X4 U35501 ( .A1(n20639), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_2), .ZN(n25585) );
NAND2_X4 U35502 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_2), .A2(n20639), .ZN(n25584) );
NAND2_X4 U35503 ( .A1(n25585), .A2(n25584), .ZN(n25586) );
NOR2_X4 U35504 ( .A1(n25587), .A2(n25586), .ZN(n25589) );
AND2_X4 U35505 ( .A1(n25587), .A2(n25586), .ZN(n25588) );
NOR2_X4 U35506 ( .A1(n25589), .A2(n25588), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_2) );
NAND2_X4 U35507 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N64), .A2(n25590), .ZN(n25593) );
OR2_X4 U35508 ( .A1(n25590), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N64), .ZN(n25591) );
NAND2_X4 U35509 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_29), .A2(n25591), .ZN(n25592) );
NAND2_X4 U35510 ( .A1(n25593), .A2(n25592), .ZN(n25599) );
OR2_X4 U35511 ( .A1(n20032), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_30), .ZN(n25595) );
NAND2_X4 U35512 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_30), .A2(n20032), .ZN(n25594) );
NAND2_X4 U35513 ( .A1(n25595), .A2(n25594), .ZN(n25596) );
NOR2_X4 U35514 ( .A1(n25599), .A2(n25596), .ZN(n25598) );
AND2_X4 U35515 ( .A1(n25599), .A2(n25596), .ZN(n25597) );
NOR2_X4 U35516 ( .A1(n25598), .A2(n25597), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_30) );
NAND2_X4 U35517 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N65), .A2(n25599), .ZN(n25602) );
OR2_X4 U35518 ( .A1(n25599), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N65), .ZN(n25600) );
NAND2_X4 U35519 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_30), .A2(n25600), .ZN(n25601) );
NAND2_X4 U35520 ( .A1(n25602), .A2(n25601), .ZN(n25608) );
OR2_X4 U35521 ( .A1(n20027), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_31), .ZN(n25604) );
NAND2_X4 U35522 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_31), .A2(n20027), .ZN(n25603) );
NAND2_X4 U35523 ( .A1(n25604), .A2(n25603), .ZN(n25605) );
NOR2_X4 U35524 ( .A1(n25608), .A2(n25605), .ZN(n25607) );
AND2_X4 U35525 ( .A1(n25608), .A2(n25605), .ZN(n25606) );
NOR2_X4 U35526 ( .A1(n25607), .A2(n25606), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_31) );
NAND2_X4 U35527 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N66), .A2(n25608), .ZN(n25611) );
OR2_X4 U35528 ( .A1(n25608), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N66), .ZN(n25609) );
NAND2_X4 U35529 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_31), .A2(n25609), .ZN(n25610) );
NAND2_X4 U35530 ( .A1(n25611), .A2(n25610), .ZN(n25619) );
OR2_X4 U35531 ( .A1(n20024), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_32), .ZN(n25613) );
NAND2_X4 U35532 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_32), .A2(n20024), .ZN(n25612) );
NAND2_X4 U35533 ( .A1(n25613), .A2(n25612), .ZN(n25614) );
NOR2_X4 U35534 ( .A1(n25619), .A2(n25614), .ZN(n25616) );
AND2_X4 U35535 ( .A1(n25619), .A2(n25614), .ZN(n25615) );
NOR2_X4 U35536 ( .A1(n25616), .A2(n25615), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_32) );
OR2_X4 U35537 ( .A1(n20025), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_33), .ZN(n25618) );
NAND2_X4 U35538 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_33), .A2(n20025), .ZN(n25617) );
NAND2_X4 U35539 ( .A1(n25618), .A2(n25617), .ZN(n25623) );
NAND2_X4 U35540 ( .A1(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N67), .A2(n25619), .ZN(n25622) );
OR2_X4 U35541 ( .A1(n25619), .A2(dp_cluster_0_ex_block_i_gen_multdiv_fast_multdiv_i_N67), .ZN(n25620) );
NAND2_X4 U35542 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_32), .A2(n25620), .ZN(n25621) );
NAND2_X4 U35543 ( .A1(n25622), .A2(n25621), .ZN(n25624) );
NOR2_X4 U35544 ( .A1(n25623), .A2(n25624), .ZN(n25626) );
AND2_X4 U35545 ( .A1(n25624), .A2(n25623), .ZN(n25625) );
NOR2_X4 U35546 ( .A1(n25626), .A2(n25625), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_33) );
OR2_X4 U35547 ( .A1(n20585), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_3), .ZN(n25628) );
NAND2_X4 U35548 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_3), .A2(n20585), .ZN(n25627) );
NAND2_X4 U35549 ( .A1(n25628), .A2(n25627), .ZN(n25629) );
NOR2_X4 U35550 ( .A1(n25630), .A2(n25629), .ZN(n25632) );
AND2_X4 U35551 ( .A1(n25630), .A2(n25629), .ZN(n25631) );
NOR2_X4 U35552 ( .A1(n25632), .A2(n25631), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_3) );
OR2_X4 U35553 ( .A1(n20546), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_4), .ZN(n25634) );
NAND2_X4 U35554 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_4), .A2(n20546), .ZN(n25633) );
NAND2_X4 U35555 ( .A1(n25634), .A2(n25633), .ZN(n25635) );
NOR2_X4 U35556 ( .A1(n25636), .A2(n25635), .ZN(n25638) );
AND2_X4 U35557 ( .A1(n25636), .A2(n25635), .ZN(n25637) );
NOR2_X4 U35558 ( .A1(n25638), .A2(n25637), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_4) );
OR2_X4 U35559 ( .A1(n20508), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_5), .ZN(n25640) );
NAND2_X4 U35560 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_5), .A2(n20508), .ZN(n25639) );
NAND2_X4 U35561 ( .A1(n25640), .A2(n25639), .ZN(n25641) );
NOR2_X4 U35562 ( .A1(n25642), .A2(n25641), .ZN(n25644) );
AND2_X4 U35563 ( .A1(n25642), .A2(n25641), .ZN(n25643) );
NOR2_X4 U35564 ( .A1(n25644), .A2(n25643), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_5) );
OR2_X4 U35565 ( .A1(n20470), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_6), .ZN(n25646) );
NAND2_X4 U35566 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_6), .A2(n20470), .ZN(n25645) );
NAND2_X4 U35567 ( .A1(n25646), .A2(n25645), .ZN(n25647) );
NOR2_X4 U35568 ( .A1(n25648), .A2(n25647), .ZN(n25650) );
AND2_X4 U35569 ( .A1(n25648), .A2(n25647), .ZN(n25649) );
NOR2_X4 U35570 ( .A1(n25650), .A2(n25649), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_6) );
OR2_X4 U35571 ( .A1(n20432), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_7), .ZN(n25652) );
NAND2_X4 U35572 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_7), .A2(n20432), .ZN(n25651) );
NAND2_X4 U35573 ( .A1(n25652), .A2(n25651), .ZN(n25653) );
NOR2_X4 U35574 ( .A1(n25654), .A2(n25653), .ZN(n25656) );
AND2_X4 U35575 ( .A1(n25654), .A2(n25653), .ZN(n25655) );
NOR2_X4 U35576 ( .A1(n25656), .A2(n25655), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_7) );
OR2_X4 U35577 ( .A1(n20395), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_8), .ZN(n25658) );
NAND2_X4 U35578 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_8), .A2(n20395), .ZN(n25657) );
NAND2_X4 U35579 ( .A1(n25658), .A2(n25657), .ZN(n25659) );
NOR2_X4 U35580 ( .A1(n25660), .A2(n25659), .ZN(n25662) );
AND2_X4 U35581 ( .A1(n25660), .A2(n25659), .ZN(n25661) );
NOR2_X4 U35582 ( .A1(n25662), .A2(n25661), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_8) );
OR2_X4 U35583 ( .A1(n20358), .A2(ex_block_i_gen_multdiv_fast_multdiv_i_accum_9), .ZN(n25664) );
NAND2_X4 U35584 ( .A1(ex_block_i_gen_multdiv_fast_multdiv_i_accum_9), .A2(n20358), .ZN(n25663) );
NAND2_X4 U35585 ( .A1(n25664), .A2(n25663), .ZN(n25665) );
NOR2_X4 U35586 ( .A1(n25666), .A2(n25665), .ZN(n25668) );
AND2_X4 U35587 ( .A1(n25666), .A2(n25665), .ZN(n25667) );
NOR2_X4 U35588 ( .A1(n25668), .A2(n25667), .ZN(ex_block_i_gen_multdiv_fast_multdiv_i_mac_res_signed_9) );
INV_X1 U35589 ( .A(n15965), .ZN(n10550) );
INV_X1 U35590 ( .A(n15964), .ZN(n10552) );
INV_X1 U35591 ( .A(n15963), .ZN(n10554) );
INV_X1 U35592 ( .A(n15962), .ZN(n10556) );
INV_X1 U35593 ( .A(n15961), .ZN(n10558) );
INV_X1 U35594 ( .A(n15960), .ZN(n10560) );
INV_X1 U35595 ( .A(n15959), .ZN(n10562) );
INV_X1 U35596 ( .A(n15958), .ZN(n10564) );
INV_X1 U35597 ( .A(n15957), .ZN(n10566) );
INV_X1 U35598 ( .A(n15956), .ZN(n10568) );
INV_X1 U35599 ( .A(n15955), .ZN(n10570) );
INV_X1 U35600 ( .A(n15954), .ZN(n10572) );
INV_X1 U35601 ( .A(n15953), .ZN(n10574) );
INV_X1 U35602 ( .A(n15952), .ZN(n10576) );
INV_X1 U35603 ( .A(n15951), .ZN(n10578) );
INV_X1 U35604 ( .A(n15950), .ZN(n10580) );
INV_X1 U35605 ( .A(n15949), .ZN(n10582) );
INV_X1 U35606 ( .A(n15948), .ZN(n10584) );
INV_X1 U35607 ( .A(n15947), .ZN(n10586) );
INV_X1 U35608 ( .A(n15946), .ZN(n10588) );
INV_X1 U35609 ( .A(n15945), .ZN(n10590) );
INV_X1 U35610 ( .A(n15944), .ZN(n10592) );
INV_X1 U35611 ( .A(n15943), .ZN(n10594) );
INV_X1 U35612 ( .A(n15942), .ZN(n10596) );
INV_X1 U35613 ( .A(n15941), .ZN(n10598) );
INV_X1 U35614 ( .A(n15940), .ZN(n10600) );
INV_X1 U35615 ( .A(n15939), .ZN(n10602) );
INV_X1 U35616 ( .A(n15938), .ZN(n10604) );
INV_X1 U35617 ( .A(n16126), .ZN(n10606) );
INV_X1 U35618 ( .A(n15937), .ZN(n10608) );
INV_X1 U35619 ( .A(crash_dump_o_5_), .ZN(n10610) );
INV_X1 U35620 ( .A(n15978), .ZN(n10612) );
INV_X1 U35621 ( .A(cs_registers_i_mhpmcounter_0__63_), .ZN(n10613) );
INV_X1 U35622 ( .A(crash_dump_o_30_), .ZN(n10615) );
INV_X1 U35623 ( .A(crash_dump_o_21_), .ZN(n10617) );
INV_X1 U35624 ( .A(crash_dump_o_29_), .ZN(n10621) );
INV_X1 U35625 ( .A(crash_dump_o_125_), .ZN(n10622) );
INV_X1 U35626 ( .A(crash_dump_o_93_), .ZN(n10623) );
INV_X1 U35627 ( .A(cs_registers_i_mhpmcounter_0__29_), .ZN(n10625) );
INV_X1 U35628 ( .A(cs_registers_i_mhpmcounter_0__61_), .ZN(n10626) );
INV_X1 U35629 ( .A(cs_registers_i_mhpmcounter_2__63_), .ZN(n10627) );
INV_X1 U35630 ( .A(cs_registers_i_mhpmcounter_2__62_), .ZN(n10628) );
INV_X1 U35631 ( .A(cs_registers_i_mhpmcounter_2__61_), .ZN(n10629) );
INV_X1 U35632 ( .A(crash_dump_o_28_), .ZN(n10631) );
INV_X1 U35633 ( .A(crash_dump_o_124_), .ZN(n10632) );
INV_X1 U35634 ( .A(crash_dump_o_92_), .ZN(n10633) );
INV_X1 U35635 ( .A(cs_registers_i_mhpmcounter_0__28_), .ZN(n10635) );
INV_X1 U35636 ( .A(cs_registers_i_mhpmcounter_0__60_), .ZN(n10636) );
INV_X1 U35637 ( .A(cs_registers_i_mhpmcounter_2__28_), .ZN(n10637) );
INV_X1 U35638 ( .A(crash_dump_o_1_), .ZN(n10644) );
INV_X1 U35639 ( .A(instr_fetch_err_plus2), .ZN(n15928) );
INV_X1 U35640 ( .A(crash_dump_o_17_), .ZN(n10646) );
INV_X1 U35641 ( .A(crash_dump_o_113_), .ZN(n10647) );
INV_X1 U35642 ( .A(crash_dump_o_81_), .ZN(n10648) );
INV_X1 U35643 ( .A(cs_registers_i_mhpmcounter_0__17_), .ZN(n10650) );
INV_X1 U35644 ( .A(cs_registers_i_mhpmcounter_0__49_), .ZN(n10651) );
INV_X1 U35645 ( .A(cs_registers_i_mhpmcounter_2__17_), .ZN(n10652) );
INV_X1 U35646 ( .A(cs_registers_i_mhpmcounter_2__49_), .ZN(n10653) );
INV_X1 U35647 ( .A(n16029), .ZN(n10654) );
INV_X1 U35648 ( .A(n16196), .ZN(n10655) );
INV_X1 U35649 ( .A(crash_dump_o_2_), .ZN(n10661) );
INV_X1 U35650 ( .A(crash_dump_o_98_), .ZN(n10662) );
INV_X1 U35651 ( .A(crash_dump_o_66_), .ZN(n10663) );
INV_X1 U35652 ( .A(cs_registers_i_mhpmcounter_0__0_), .ZN(n10665) );
INV_X1 U35653 ( .A(cs_registers_i_mhpmcounter_0__1_), .ZN(n10666) );
INV_X1 U35654 ( .A(cs_registers_i_mhpmcounter_0__2_), .ZN(n10667) );
INV_X1 U35655 ( .A(crash_dump_o_3_), .ZN(n10669) );
INV_X1 U35656 ( .A(crash_dump_o_99_), .ZN(n10670) );
INV_X1 U35657 ( .A(crash_dump_o_67_), .ZN(n10671) );
INV_X1 U35658 ( .A(cs_registers_i_mhpmcounter_0__35_), .ZN(n10673) );
INV_X1 U35659 ( .A(cs_registers_i_mhpmcounter_2__35_), .ZN(n10674) );
INV_X1 U35660 ( .A(cs_registers_i_mhpmcounter_2__3_), .ZN(n10675) );
INV_X1 U35661 ( .A(n16050), .ZN(n10677) );
INV_X1 U35662 ( .A(crash_dump_o_7_), .ZN(n10679) );
INV_X1 U35663 ( .A(crash_dump_o_103_), .ZN(n10680) );
INV_X1 U35664 ( .A(crash_dump_o_71_), .ZN(n10681) );
INV_X1 U35665 ( .A(cs_registers_i_mhpmcounter_0__39_), .ZN(n10683) );
INV_X1 U35666 ( .A(cs_registers_i_mhpmcounter_0__7_), .ZN(n10684) );
INV_X1 U35667 ( .A(cs_registers_i_mhpmcounter_2__39_), .ZN(n10685) );
INV_X1 U35668 ( .A(cs_registers_i_mhpmcounter_2__7_), .ZN(n10686) );
INV_X1 U35669 ( .A(n15977), .ZN(n10692) );
INV_X1 U35670 ( .A(cs_registers_i_mhpmcounter_0__36_), .ZN(n10693) );
INV_X1 U35671 ( .A(cs_registers_i_mhpmcounter_0__4_), .ZN(n10694) );
INV_X1 U35672 ( .A(cs_registers_i_mhpmcounter_2__36_), .ZN(n10695) );
INV_X1 U35673 ( .A(cs_registers_i_mhpmcounter_2__4_), .ZN(n10696) );
INV_X1 U35674 ( .A(crash_dump_o_4_), .ZN(n10698) );
INV_X1 U35675 ( .A(crash_dump_o_100_), .ZN(n10704) );
INV_X1 U35676 ( .A(crash_dump_o_68_), .ZN(n10705) );
INV_X1 U35677 ( .A(cs_registers_i_mhpmcounter_0__38_), .ZN(n10706) );
INV_X1 U35678 ( .A(cs_registers_i_mhpmcounter_0__6_), .ZN(n10707) );
INV_X1 U35679 ( .A(cs_registers_i_mhpmcounter_2__38_), .ZN(n10708) );
INV_X1 U35680 ( .A(cs_registers_i_mhpmcounter_2__6_), .ZN(n10709) );
INV_X1 U35681 ( .A(crash_dump_o_6_), .ZN(n10711) );
INV_X1 U35682 ( .A(crash_dump_o_102_), .ZN(n10717) );
INV_X1 U35683 ( .A(crash_dump_o_70_), .ZN(n10718) );
INV_X1 U35684 ( .A(cs_registers_i_mhpmcounter_0__40_), .ZN(n10719) );
INV_X1 U35685 ( .A(cs_registers_i_mhpmcounter_0__8_), .ZN(n10720) );
INV_X1 U35686 ( .A(cs_registers_i_mhpmcounter_2__40_), .ZN(n10721) );
INV_X1 U35687 ( .A(cs_registers_i_mhpmcounter_2__8_), .ZN(n10722) );
INV_X1 U35688 ( .A(n16023), .ZN(n10723) );
INV_X1 U35689 ( .A(crash_dump_o_8_), .ZN(n10725) );
INV_X1 U35690 ( .A(crash_dump_o_104_), .ZN(n10731) );
INV_X1 U35691 ( .A(crash_dump_o_72_), .ZN(n10732) );
INV_X1 U35692 ( .A(cs_registers_i_mhpmcounter_0__41_), .ZN(n10733) );
INV_X1 U35693 ( .A(cs_registers_i_mhpmcounter_0__9_), .ZN(n10734) );
INV_X1 U35694 ( .A(cs_registers_i_mhpmcounter_2__41_), .ZN(n10735) );
INV_X1 U35695 ( .A(cs_registers_i_mhpmcounter_2__9_), .ZN(n10736) );
INV_X1 U35696 ( .A(n16039), .ZN(n10737) );
INV_X1 U35697 ( .A(crash_dump_o_9_), .ZN(n10739) );
INV_X1 U35698 ( .A(crash_dump_o_105_), .ZN(n10745) );
INV_X1 U35699 ( .A(crash_dump_o_73_), .ZN(n10746) );
INV_X1 U35700 ( .A(cs_registers_i_mhpmcounter_0__10_), .ZN(n10747) );
INV_X1 U35701 ( .A(cs_registers_i_mhpmcounter_0__42_), .ZN(n10748) );
INV_X1 U35702 ( .A(cs_registers_i_mhpmcounter_2__10_), .ZN(n10749) );
INV_X1 U35703 ( .A(cs_registers_i_mhpmcounter_2__42_), .ZN(n10750) );
INV_X1 U35704 ( .A(n16024), .ZN(n10751) );
INV_X1 U35705 ( .A(crash_dump_o_10_), .ZN(n10753) );
INV_X1 U35706 ( .A(crash_dump_o_106_), .ZN(n10759) );
INV_X1 U35707 ( .A(crash_dump_o_74_), .ZN(n10760) );
INV_X1 U35708 ( .A(cs_registers_i_mhpmcounter_0__11_), .ZN(n10761) );
INV_X1 U35709 ( .A(cs_registers_i_mhpmcounter_0__43_), .ZN(n10762) );
INV_X1 U35710 ( .A(cs_registers_i_mhpmcounter_2__11_), .ZN(n10763) );
INV_X1 U35711 ( .A(cs_registers_i_mhpmcounter_2__43_), .ZN(n10764) );
INV_X1 U35712 ( .A(n16133), .ZN(n10766) );
INV_X1 U35713 ( .A(crash_dump_o_12_), .ZN(n10768) );
INV_X1 U35714 ( .A(crash_dump_o_108_), .ZN(n10769) );
INV_X1 U35715 ( .A(crash_dump_o_76_), .ZN(n10770) );
INV_X1 U35716 ( .A(cs_registers_i_mhpmcounter_0__12_), .ZN(n10772) );
INV_X1 U35717 ( .A(cs_registers_i_mhpmcounter_0__44_), .ZN(n10773) );
INV_X1 U35718 ( .A(cs_registers_i_mhpmcounter_2__12_), .ZN(n10774) );
INV_X1 U35719 ( .A(cs_registers_i_mhpmcounter_2__44_), .ZN(n10775) );
INV_X1 U35720 ( .A(n16025), .ZN(n10776) );
INV_X1 U35721 ( .A(priv_mode_id_1), .ZN(n15817) );
INV_X1 U35722 ( .A(cs_registers_i_mhpmcounter_0__13_), .ZN(n10782) );
INV_X1 U35723 ( .A(cs_registers_i_mhpmcounter_0__45_), .ZN(n10783) );
INV_X1 U35724 ( .A(cs_registers_i_mhpmcounter_2__13_), .ZN(n10784) );
INV_X1 U35725 ( .A(cs_registers_i_mhpmcounter_2__45_), .ZN(n10785) );
INV_X1 U35726 ( .A(crash_dump_o_13_), .ZN(n10787) );
INV_X1 U35727 ( .A(crash_dump_o_109_), .ZN(n10788) );
INV_X1 U35728 ( .A(crash_dump_o_77_), .ZN(n10789) );
INV_X1 U35729 ( .A(n16026), .ZN(n10790) );
INV_X1 U35730 ( .A(cs_registers_i_mhpmcounter_0__14_), .ZN(n10797) );
INV_X1 U35731 ( .A(cs_registers_i_mhpmcounter_0__46_), .ZN(n10798) );
INV_X1 U35732 ( .A(cs_registers_i_mhpmcounter_2__14_), .ZN(n10799) );
INV_X1 U35733 ( .A(cs_registers_i_mhpmcounter_2__46_), .ZN(n10800) );
INV_X1 U35734 ( .A(crash_dump_o_14_), .ZN(n10802) );
INV_X1 U35735 ( .A(crash_dump_o_110_), .ZN(n10803) );
INV_X1 U35736 ( .A(crash_dump_o_78_), .ZN(n10804) );
INV_X1 U35737 ( .A(n16027), .ZN(n10805) );
INV_X1 U35738 ( .A(cs_registers_i_mhpmcounter_0__15_), .ZN(n10811) );
INV_X1 U35739 ( .A(cs_registers_i_mhpmcounter_0__47_), .ZN(n10812) );
INV_X1 U35740 ( .A(cs_registers_i_mhpmcounter_2__15_), .ZN(n10813) );
INV_X1 U35741 ( .A(cs_registers_i_mhpmcounter_2__47_), .ZN(n10814) );
INV_X1 U35742 ( .A(crash_dump_o_15_), .ZN(n10816) );
INV_X1 U35743 ( .A(crash_dump_o_111_), .ZN(n10817) );
INV_X1 U35744 ( .A(crash_dump_o_79_), .ZN(n10818) );
INV_X1 U35745 ( .A(n16028), .ZN(n10819) );
INV_X1 U35746 ( .A(n16043), .ZN(n10820) );
INV_X1 U35747 ( .A(cs_registers_i_mhpmcounter_0__16_), .ZN(n10826) );
INV_X1 U35748 ( .A(cs_registers_i_mhpmcounter_0__48_), .ZN(n10827) );
INV_X1 U35749 ( .A(cs_registers_i_mhpmcounter_2__16_), .ZN(n10828) );
INV_X1 U35750 ( .A(cs_registers_i_mhpmcounter_2__48_), .ZN(n10829) );
INV_X1 U35751 ( .A(crash_dump_o_16_), .ZN(n10831) );
INV_X1 U35752 ( .A(crash_dump_o_112_), .ZN(n10832) );
INV_X1 U35753 ( .A(crash_dump_o_80_), .ZN(n10833) );
INV_X1 U35754 ( .A(n16017), .ZN(n10839) );
INV_X1 U35755 ( .A(cs_registers_i_mhpmcounter_0__18_), .ZN(n10841) );
INV_X1 U35756 ( .A(cs_registers_i_mhpmcounter_0__50_), .ZN(n10842) );
INV_X1 U35757 ( .A(cs_registers_i_mhpmcounter_2__18_), .ZN(n10843) );
INV_X1 U35758 ( .A(cs_registers_i_mhpmcounter_2__50_), .ZN(n10844) );
INV_X1 U35759 ( .A(crash_dump_o_18_), .ZN(n10846) );
INV_X1 U35760 ( .A(crash_dump_o_114_), .ZN(n10847) );
INV_X1 U35761 ( .A(crash_dump_o_82_), .ZN(n10848) );
INV_X1 U35762 ( .A(n16030), .ZN(n10849) );
INV_X1 U35763 ( .A(n16049), .ZN(n10855) );
INV_X1 U35764 ( .A(n16006), .ZN(n10856) );
INV_X1 U35765 ( .A(cs_registers_i_mhpmcounter_0__19_), .ZN(n10858) );
INV_X1 U35766 ( .A(cs_registers_i_mhpmcounter_0__51_), .ZN(n10859) );
INV_X1 U35767 ( .A(cs_registers_i_mhpmcounter_2__19_), .ZN(n10860) );
INV_X1 U35768 ( .A(cs_registers_i_mhpmcounter_2__51_), .ZN(n10861) );
INV_X1 U35769 ( .A(crash_dump_o_19_), .ZN(n10863) );
INV_X1 U35770 ( .A(crash_dump_o_115_), .ZN(n10864) );
INV_X1 U35771 ( .A(crash_dump_o_83_), .ZN(n10865) );
INV_X1 U35772 ( .A(n16031), .ZN(n10866) );
INV_X1 U35773 ( .A(n16012), .ZN(n10871) );
INV_X1 U35774 ( .A(cs_registers_i_mhpmcounter_0__20_), .ZN(n10873) );
INV_X1 U35775 ( .A(cs_registers_i_mhpmcounter_0__52_), .ZN(n10874) );
INV_X1 U35776 ( .A(cs_registers_i_mhpmcounter_2__20_), .ZN(n10875) );
INV_X1 U35777 ( .A(cs_registers_i_mhpmcounter_2__52_), .ZN(n10876) );
INV_X1 U35778 ( .A(crash_dump_o_20_), .ZN(n10878) );
INV_X1 U35779 ( .A(crash_dump_o_116_), .ZN(n10879) );
INV_X1 U35780 ( .A(crash_dump_o_84_), .ZN(n10880) );
INV_X1 U35781 ( .A(n16013), .ZN(n10886) );
INV_X1 U35782 ( .A(cs_registers_i_mhpmcounter_0__22_), .ZN(n10888) );
INV_X1 U35783 ( .A(cs_registers_i_mhpmcounter_0__54_), .ZN(n10889) );
INV_X1 U35784 ( .A(cs_registers_i_mhpmcounter_2__22_), .ZN(n10890) );
INV_X1 U35785 ( .A(cs_registers_i_mhpmcounter_2__54_), .ZN(n10891) );
INV_X1 U35786 ( .A(crash_dump_o_22_), .ZN(n10893) );
INV_X1 U35787 ( .A(crash_dump_o_118_), .ZN(n10894) );
INV_X1 U35788 ( .A(crash_dump_o_86_), .ZN(n10895) );
INV_X1 U35789 ( .A(n16033), .ZN(n10896) );
INV_X1 U35790 ( .A(n16003), .ZN(n10901) );
INV_X1 U35791 ( .A(cs_registers_i_mhpmcounter_0__23_), .ZN(n10903) );
INV_X1 U35792 ( .A(cs_registers_i_mhpmcounter_0__55_), .ZN(n10904) );
INV_X1 U35793 ( .A(cs_registers_i_mhpmcounter_2__23_), .ZN(n10905) );
INV_X1 U35794 ( .A(cs_registers_i_mhpmcounter_2__55_), .ZN(n10906) );
INV_X1 U35795 ( .A(crash_dump_o_23_), .ZN(n10908) );
INV_X1 U35796 ( .A(crash_dump_o_119_), .ZN(n10909) );
INV_X1 U35797 ( .A(crash_dump_o_87_), .ZN(n10910) );
INV_X1 U35798 ( .A(n16034), .ZN(n10911) );
INV_X1 U35799 ( .A(n16010), .ZN(n10916) );
INV_X1 U35800 ( .A(cs_registers_i_mhpmcounter_0__24_), .ZN(n10918) );
INV_X1 U35801 ( .A(cs_registers_i_mhpmcounter_0__56_), .ZN(n10919) );
INV_X1 U35802 ( .A(cs_registers_i_mhpmcounter_2__24_), .ZN(n10920) );
INV_X1 U35803 ( .A(cs_registers_i_mhpmcounter_2__56_), .ZN(n10921) );
INV_X1 U35804 ( .A(crash_dump_o_24_), .ZN(n10923) );
INV_X1 U35805 ( .A(crash_dump_o_120_), .ZN(n10924) );
INV_X1 U35806 ( .A(crash_dump_o_88_), .ZN(n10925) );
INV_X1 U35807 ( .A(n16035), .ZN(n10926) );
INV_X1 U35808 ( .A(n16009), .ZN(n10931) );
INV_X1 U35809 ( .A(cs_registers_i_mhpmcounter_0__25_), .ZN(n10933) );
INV_X1 U35810 ( .A(cs_registers_i_mhpmcounter_0__57_), .ZN(n10934) );
INV_X1 U35811 ( .A(cs_registers_i_mhpmcounter_2__25_), .ZN(n10935) );
INV_X1 U35812 ( .A(cs_registers_i_mhpmcounter_2__57_), .ZN(n10936) );
INV_X1 U35813 ( .A(crash_dump_o_25_), .ZN(n10938) );
INV_X1 U35814 ( .A(crash_dump_o_121_), .ZN(n10939) );
INV_X1 U35815 ( .A(crash_dump_o_89_), .ZN(n10940) );
INV_X1 U35816 ( .A(n16000), .ZN(n10946) );
INV_X1 U35817 ( .A(cs_registers_i_mhpmcounter_0__26_), .ZN(n10948) );
INV_X1 U35818 ( .A(cs_registers_i_mhpmcounter_0__58_), .ZN(n10949) );
INV_X1 U35819 ( .A(cs_registers_i_mhpmcounter_2__26_), .ZN(n10950) );
INV_X1 U35820 ( .A(cs_registers_i_mhpmcounter_2__58_), .ZN(n10951) );
INV_X1 U35821 ( .A(crash_dump_o_26_), .ZN(n10953) );
INV_X1 U35822 ( .A(crash_dump_o_122_), .ZN(n10954) );
INV_X1 U35823 ( .A(crash_dump_o_90_), .ZN(n10955) );
INV_X1 U35824 ( .A(n16036), .ZN(n10956) );
INV_X1 U35825 ( .A(n16001), .ZN(n10961) );
INV_X1 U35826 ( .A(cs_registers_i_mhpmcounter_0__27_), .ZN(n10963) );
INV_X1 U35827 ( .A(cs_registers_i_mhpmcounter_0__59_), .ZN(n10964) );
INV_X1 U35828 ( .A(cs_registers_i_mhpmcounter_2__27_), .ZN(n10965) );
INV_X1 U35829 ( .A(cs_registers_i_mhpmcounter_2__59_), .ZN(n10966) );
INV_X1 U35830 ( .A(crash_dump_o_27_), .ZN(n10968) );
INV_X1 U35831 ( .A(crash_dump_o_123_), .ZN(n10969) );
INV_X1 U35832 ( .A(crash_dump_o_91_), .ZN(n10970) );
INV_X1 U35833 ( .A(n16004), .ZN(n10976) );
INV_X1 U35834 ( .A(crash_dump_o_11_), .ZN(n10979) );
INV_X1 U35835 ( .A(crash_dump_o_31_), .ZN(n10981) );
INV_X1 U35836 ( .A(crash_dump_o_0_), .ZN(n11008) );
INV_X1 U35837 ( .A(nmi_mode), .ZN(n15919) );
INV_X1 U35838 ( .A(n15798), .ZN(n11515) );
INV_X1 U35839 ( .A(n16032), .ZN(n11019) );
INV_X1 U35840 ( .A(n16037), .ZN(n11020) );
INV_X1 U35841 ( .A(n16038), .ZN(n11021) );
INV_X1 U35842 ( .A(n16040), .ZN(n11022) );
INV_X1 U35843 ( .A(crash_dump_o_33_), .ZN(n11031) );
INV_X1 U35844 ( .A(crash_dump_o_34_), .ZN(n11032) );
INV_X1 U35845 ( .A(crash_dump_o_35_), .ZN(n11033) );
INV_X1 U35846 ( .A(crash_dump_o_36_), .ZN(n11034) );
INV_X1 U35847 ( .A(crash_dump_o_38_), .ZN(n11036) );
INV_X1 U35848 ( .A(crash_dump_o_39_), .ZN(n11037) );
INV_X1 U35849 ( .A(crash_dump_o_40_), .ZN(n11038) );
INV_X1 U35850 ( .A(crash_dump_o_41_), .ZN(n11039) );
INV_X1 U35851 ( .A(crash_dump_o_42_), .ZN(n11040) );
INV_X1 U35852 ( .A(crash_dump_o_44_), .ZN(n11042) );
INV_X1 U35853 ( .A(crash_dump_o_45_), .ZN(n11043) );
INV_X1 U35854 ( .A(crash_dump_o_46_), .ZN(n11044) );
INV_X1 U35855 ( .A(crash_dump_o_47_), .ZN(n11045) );
INV_X1 U35856 ( .A(crash_dump_o_48_), .ZN(n11046) );
INV_X1 U35857 ( .A(crash_dump_o_49_), .ZN(n11047) );
INV_X1 U35858 ( .A(crash_dump_o_50_), .ZN(n11048) );
INV_X1 U35859 ( .A(crash_dump_o_51_), .ZN(n11049) );
INV_X1 U35860 ( .A(crash_dump_o_52_), .ZN(n11050) );
INV_X1 U35861 ( .A(crash_dump_o_53_), .ZN(n11051) );
INV_X1 U35862 ( .A(crash_dump_o_54_), .ZN(n11052) );
INV_X1 U35863 ( .A(crash_dump_o_55_), .ZN(n11053) );
INV_X1 U35864 ( .A(crash_dump_o_56_), .ZN(n11054) );
INV_X1 U35865 ( .A(crash_dump_o_57_), .ZN(n11055) );
INV_X1 U35866 ( .A(crash_dump_o_58_), .ZN(n11056) );
INV_X1 U35867 ( .A(crash_dump_o_59_), .ZN(n11057) );
INV_X1 U35868 ( .A(crash_dump_o_60_), .ZN(n11058) );
INV_X1 U35869 ( .A(crash_dump_o_61_), .ZN(n11492) );
INV_X1 U35870 ( .A(crash_dump_o_62_), .ZN(n11059) );
INV_X1 U35871 ( .A(crash_dump_o_63_), .ZN(n11060) );
INV_X1 U35872 ( .A(crash_dump_o_32_), .ZN(n11061) );
INV_X1 U35873 ( .A(n15923), .ZN(n11062) );
INV_X1 U35874 ( .A(n16115), .ZN(n11064) );
INV_X1 U35875 ( .A(n16073), .ZN(n11073) );
INV_X1 U35876 ( .A(n16072), .ZN(n11074) );
INV_X1 U35877 ( .A(n16071), .ZN(n11075) );
INV_X1 U35878 ( .A(n16070), .ZN(n11076) );
INV_X1 U35879 ( .A(n16069), .ZN(n11077) );
INV_X1 U35880 ( .A(n16068), .ZN(n11078) );
INV_X1 U35881 ( .A(n16067), .ZN(n11079) );
INV_X1 U35882 ( .A(n16066), .ZN(n11080) );
INV_X1 U35883 ( .A(n16065), .ZN(n11081) );
INV_X1 U35884 ( .A(n16064), .ZN(n11082) );
INV_X1 U35885 ( .A(n16063), .ZN(n11083) );
INV_X1 U35886 ( .A(n16062), .ZN(n11084) );
INV_X1 U35887 ( .A(n16061), .ZN(n11085) );
INV_X1 U35888 ( .A(n16060), .ZN(n11086) );
INV_X1 U35889 ( .A(n16059), .ZN(n11087) );
INV_X1 U35890 ( .A(n16058), .ZN(n11088) );
INV_X1 U35891 ( .A(n15911), .ZN(n11090) );
INV_X1 U35892 ( .A(n15822), .ZN(n11091) );
INV_X1 U35893 ( .A(cs_registers_i_mhpmcounter_0__21_), .ZN(n11114) );
INV_X1 U35894 ( .A(cs_registers_i_mhpmcounter_0__30_), .ZN(n11115) );
INV_X1 U35895 ( .A(cs_registers_i_mhpmcounter_0__32_), .ZN(n11116) );
INV_X1 U35896 ( .A(cs_registers_i_mhpmcounter_0__33_), .ZN(n11117) );
INV_X1 U35897 ( .A(cs_registers_i_mhpmcounter_0__34_), .ZN(n11118) );
INV_X1 U35898 ( .A(cs_registers_i_mhpmcounter_0__37_), .ZN(n11119) );
INV_X1 U35899 ( .A(cs_registers_i_mhpmcounter_0__53_), .ZN(n11120) );
INV_X1 U35900 ( .A(cs_registers_i_mhpmcounter_0__5_), .ZN(n11121) );
INV_X1 U35901 ( .A(cs_registers_i_mhpmcounter_2__1_), .ZN(n11122) );
INV_X1 U35902 ( .A(cs_registers_i_mhpmcounter_2__21_), .ZN(n11123) );
INV_X1 U35903 ( .A(cs_registers_i_mhpmcounter_2__2_), .ZN(n11124) );
INV_X1 U35904 ( .A(cs_registers_i_mhpmcounter_2__30_), .ZN(n11125) );
INV_X1 U35905 ( .A(cs_registers_i_mhpmcounter_2__31_), .ZN(n11126) );
INV_X1 U35906 ( .A(cs_registers_i_mhpmcounter_2__32_), .ZN(n11127) );
INV_X1 U35907 ( .A(cs_registers_i_mhpmcounter_2__33_), .ZN(n11128) );
INV_X1 U35908 ( .A(cs_registers_i_mhpmcounter_2__34_), .ZN(n11129) );
INV_X1 U35909 ( .A(cs_registers_i_mhpmcounter_2__37_), .ZN(n11130) );
INV_X1 U35910 ( .A(cs_registers_i_mhpmcounter_2__53_), .ZN(n11131) );
INV_X1 U35911 ( .A(cs_registers_i_mhpmcounter_2__5_), .ZN(n11132) );
INV_X1 U35912 ( .A(n16015), .ZN(n11144) );
INV_X1 U35913 ( .A(n16016), .ZN(n11145) );
INV_X1 U35914 ( .A(n16127), .ZN(n11146) );
INV_X1 U35915 ( .A(n16008), .ZN(n11147) );
INV_X1 U35916 ( .A(n16011), .ZN(n11148) );
INV_X1 U35917 ( .A(n16125), .ZN(n11500) );
INV_X1 U35918 ( .A(n15931), .ZN(n11153) );
INV_X1 U35919 ( .A(n15930), .ZN(n11154) );
INV_X1 U35920 ( .A(n15906), .ZN(n11156) );
INV_X1 U35921 ( .A(n15905), .ZN(n11157) );
INV_X1 U35922 ( .A(n15904), .ZN(n11158) );
INV_X1 U35923 ( .A(n15903), .ZN(n11159) );
INV_X1 U35924 ( .A(n15902), .ZN(n11160) );
INV_X1 U35925 ( .A(n15901), .ZN(n11161) );
INV_X1 U35926 ( .A(n15900), .ZN(n11162) );
INV_X1 U35927 ( .A(n15899), .ZN(n11163) );
INV_X1 U35928 ( .A(n15898), .ZN(n11164) );
INV_X1 U35929 ( .A(n15886), .ZN(n11165) );
INV_X1 U35930 ( .A(n16194), .ZN(n11217) );
INV_X1 U35931 ( .A(n16193), .ZN(n11185) );
INV_X1 U35932 ( .A(n15875), .ZN(n11166) );
INV_X1 U35933 ( .A(n15874), .ZN(n11167) );
INV_X1 U35934 ( .A(n15873), .ZN(n11168) );
INV_X1 U35935 ( .A(n15872), .ZN(n11169) );
INV_X1 U35936 ( .A(n15871), .ZN(n11170) );
INV_X1 U35937 ( .A(n15870), .ZN(n11171) );
INV_X1 U35938 ( .A(n15869), .ZN(n11172) );
INV_X1 U35939 ( .A(n15868), .ZN(n11173) );
INV_X1 U35940 ( .A(n15867), .ZN(n11174) );
INV_X1 U35941 ( .A(n15866), .ZN(n11175) );
INV_X1 U35942 ( .A(n15865), .ZN(n11176) );
INV_X1 U35943 ( .A(n15864), .ZN(n11177) );
INV_X1 U35944 ( .A(n15863), .ZN(n11178) );
INV_X1 U35945 ( .A(n15862), .ZN(n11179) );
INV_X1 U35946 ( .A(n15861), .ZN(n11180) );
INV_X1 U35947 ( .A(n15883), .ZN(n11181) );
INV_X1 U35948 ( .A(n15882), .ZN(n11182) );
INV_X1 U35949 ( .A(n15881), .ZN(n11183) );
INV_X1 U35950 ( .A(n15880), .ZN(n11184) );
INV_X1 U35951 ( .A(n15897), .ZN(n11186) );
INV_X1 U35952 ( .A(n16192), .ZN(n11187) );
INV_X1 U35953 ( .A(n16191), .ZN(n11188) );
INV_X1 U35954 ( .A(n16190), .ZN(n11189) );
INV_X1 U35955 ( .A(n16189), .ZN(n11190) );
INV_X1 U35956 ( .A(n16188), .ZN(n11191) );
INV_X1 U35957 ( .A(n16187), .ZN(n11192) );
INV_X1 U35958 ( .A(n16186), .ZN(n11193) );
INV_X1 U35959 ( .A(n16185), .ZN(n11194) );
INV_X1 U35960 ( .A(n16184), .ZN(n11195) );
INV_X1 U35961 ( .A(n16183), .ZN(n11196) );
INV_X1 U35962 ( .A(n16182), .ZN(n11197) );
INV_X1 U35963 ( .A(n16181), .ZN(n11198) );
INV_X1 U35964 ( .A(n16180), .ZN(n11199) );
INV_X1 U35965 ( .A(n16179), .ZN(n11200) );
INV_X1 U35966 ( .A(n16178), .ZN(n11201) );
INV_X1 U35967 ( .A(n16177), .ZN(n11202) );
INV_X1 U35968 ( .A(n16176), .ZN(n11203) );
INV_X1 U35969 ( .A(n16175), .ZN(n11204) );
INV_X1 U35970 ( .A(n16174), .ZN(n11205) );
INV_X1 U35971 ( .A(n16173), .ZN(n11206) );
INV_X1 U35972 ( .A(n16172), .ZN(n11207) );
INV_X1 U35973 ( .A(n16153), .ZN(n11215) );
INV_X1 U35974 ( .A(n16152), .ZN(n11208) );
INV_X1 U35975 ( .A(n16151), .ZN(n11209) );
INV_X1 U35976 ( .A(n16150), .ZN(n11210) );
INV_X1 U35977 ( .A(n16149), .ZN(n11211) );
INV_X1 U35978 ( .A(n16148), .ZN(n11212) );
INV_X1 U35979 ( .A(n16147), .ZN(n11213) );
INV_X1 U35980 ( .A(n16146), .ZN(n11214) );
INV_X1 U35981 ( .A(n15891), .ZN(n11216) );
INV_X1 U35982 ( .A(n15896), .ZN(n11218) );
INV_X1 U35983 ( .A(n16171), .ZN(n11220) );
INV_X1 U35984 ( .A(n16170), .ZN(n11221) );
INV_X1 U35985 ( .A(n16169), .ZN(n11222) );
INV_X1 U35986 ( .A(n16168), .ZN(n11231) );
INV_X1 U35987 ( .A(n16167), .ZN(n11242) );
INV_X1 U35988 ( .A(n16041), .ZN(n11244) );
INV_X1 U35989 ( .A(n16144), .ZN(n11245) );
INV_X1 U35990 ( .A(n16143), .ZN(n11246) );
INV_X1 U35991 ( .A(n16142), .ZN(n11247) );
INV_X1 U35992 ( .A(n16141), .ZN(n11248) );
INV_X1 U35993 ( .A(n16140), .ZN(n11249) );
INV_X1 U35994 ( .A(n16139), .ZN(n11250) );
INV_X1 U35995 ( .A(n16138), .ZN(n11251) );
INV_X1 U35996 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_4), .ZN(n11252) );
INV_X1 U35997 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_3), .ZN(n11253) );
INV_X1 U35998 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_2), .ZN(n11254) );
INV_X1 U35999 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_1), .ZN(n11255) );
INV_X1 U36000 ( .A(ex_block_i_gen_multdiv_fast_multdiv_i_div_counter_q_0), .ZN(n11256) );
INV_X1 U36001 ( .A(n15887), .ZN(n11289) );
INV_X1 U36002 ( .A(n16166), .ZN(n11257) );
INV_X1 U36003 ( .A(n16165), .ZN(n11258) );
INV_X1 U36004 ( .A(n16164), .ZN(n11259) );
INV_X1 U36005 ( .A(n16163), .ZN(n11262) );
INV_X1 U36006 ( .A(n16162), .ZN(n11263) );
INV_X1 U36007 ( .A(n16161), .ZN(n11264) );
INV_X1 U36008 ( .A(n16160), .ZN(n11265) );
INV_X1 U36009 ( .A(n16159), .ZN(n11266) );
INV_X1 U36010 ( .A(n16158), .ZN(n11267) );
INV_X1 U36011 ( .A(n16157), .ZN(n11274) );
INV_X1 U36012 ( .A(n16156), .ZN(n11277) );
INV_X1 U36013 ( .A(n16155), .ZN(n11278) );
INV_X1 U36014 ( .A(n16154), .ZN(n11279) );
INV_X1 U36015 ( .A(n16084), .ZN(n11281) );
INV_X1 U36016 ( .A(n16137), .ZN(n11282) );
INV_X1 U36017 ( .A(n16136), .ZN(n11285) );
INV_X1 U36018 ( .A(n16135), .ZN(n11286) );
INV_X1 U36019 ( .A(n16134), .ZN(n11287) );
INV_X1 U36020 ( .A(n15877), .ZN(n11290) );
INV_X1 U36021 ( .A(n15888), .ZN(n11291) );
INV_X1 U36022 ( .A(n16197), .ZN(n11292) );
INV_X1 U36023 ( .A(n15916), .ZN(n11293) );
INV_X1 U36024 ( .A(n16131), .ZN(n11294) );
INV_X1 U36025 ( .A(n15925), .ZN(n11295) );
INV_X1 U36026 ( .A(n16130), .ZN(n11297) );
INV_X1 U36027 ( .A(n15825), .ZN(n11296) );
INV_X1 U36028 ( .A(n16145), .ZN(n11298) );
INV_X1 U36029 ( .A(n15922), .ZN(n11299) );
INV_X1 U36030 ( .A(n15823), .ZN(n11300) );
INV_X1 U36031 ( .A(n15915), .ZN(n11516) );
INV_X1 U36032 ( .A(n15909), .ZN(n11301) );
INV_X1 U36033 ( .A(n15813), .ZN(n11498) );
INV_X1 U36034 ( .A(n15819), .ZN(n11514) );
INV_X1 U36035 ( .A(n16042), .ZN(n11302) );
INV_X1 U36036 ( .A(n15907), .ZN(n11519) );
INV_X1 U36037 ( .A(priv_mode_id_0), .ZN(n15913) );
INV_X1 U36038 ( .A(crash_dump_o_107_), .ZN(n11307) );
INV_X1 U36039 ( .A(crash_dump_o_75_), .ZN(n11308) );
INV_X1 U36040 ( .A(n15800), .ZN(n11517) );
INV_X1 U36041 ( .A(rf_waddr_wb_o_3_), .ZN(n15826) );
INV_X1 U36042 ( .A(rf_waddr_wb_o_4_), .ZN(n16082) );
INV_X1 U36043 ( .A(rf_raddr_b_o_4_), .ZN(n11311) );
INV_X1 U36044 ( .A(n15893), .ZN(n11312) );
INV_X1 U36045 ( .A(n15858), .ZN(n11313) );
INV_X1 U36046 ( .A(rf_raddr_a_o_4_), .ZN(n15885) );
INV_X1 U36047 ( .A(n15918), .ZN(n11493) );
INV_X1 U36048 ( .A(n15924), .ZN(n11316) );
INV_X1 U36049 ( .A(n15814), .ZN(n11317) );
INV_X1 U36050 ( .A(n15884), .ZN(n11318) );
INV_X1 U36051 ( .A(n15810), .ZN(n11319) );
INV_X1 U36052 ( .A(n15879), .ZN(n11320) );
INV_X1 U36053 ( .A(n15912), .ZN(n11321) );
INV_X1 U36054 ( .A(n15895), .ZN(n11501) );
INV_X1 U36055 ( .A(n15799), .ZN(n11322) );
INV_X1 U36056 ( .A(n15917), .ZN(n11504) );
INV_X1 U36057 ( .A(rf_raddr_a_o_0_), .ZN(n15890) );
INV_X1 U36058 ( .A(rf_raddr_a_o_2_), .ZN(n15889) );
INV_X1 U36059 ( .A(rf_raddr_b_o_2_), .ZN(n11323) );
INV_X1 U36060 ( .A(n15816), .ZN(n11324) );
INV_X1 U36061 ( .A(n15807), .ZN(n11325) );
INV_X1 U36062 ( .A(n15908), .ZN(n11326) );
INV_X1 U36063 ( .A(n15876), .ZN(n11502) );
INV_X1 U36064 ( .A(n15910), .ZN(n11327) );
INV_X1 U36065 ( .A(n15804), .ZN(n11503) );
INV_X1 U36066 ( .A(n15859), .ZN(n11328) );
INV_X1 U36067 ( .A(n15805), .ZN(n11329) );
INV_X1 U36068 ( .A(rf_raddr_a_o_1_), .ZN(n15809) );
INV_X1 U36069 ( .A(rf_raddr_a_o_3_), .ZN(n15806) );
INV_X1 U36070 ( .A(rf_raddr_b_o_0_), .ZN(n11330) );
INV_X1 U36071 ( .A(rf_raddr_b_o_1_), .ZN(n11331) );
INV_X1 U36072 ( .A(rf_raddr_b_o_3_), .ZN(n11332) );
INV_X1 U36073 ( .A(n15914), .ZN(n11333) );
INV_X1 U36074 ( .A(n15824), .ZN(n11334) );
INV_X1 U36075 ( .A(n15815), .ZN(n11336) );
INV_X1 U36076 ( .A(n15982), .ZN(n11338) );
INV_X1 U36077 ( .A(n16128), .ZN(n11339) );
INV_X1 U36078 ( .A(n15892), .ZN(n11340) );
INV_X1 U36079 ( .A(rf_waddr_wb_o_0_), .ZN(n16123) );
INV_X1 U36080 ( .A(rf_waddr_wb_o_1_), .ZN(n15828) );
INV_X1 U36081 ( .A(n15894), .ZN(n11345) );
INV_X1 U36082 ( .A(n15970), .ZN(n11375) );
INV_X1 U36083 ( .A(n15969), .ZN(n11380) );
INV_X1 U36084 ( .A(n15968), .ZN(n11383) );
INV_X1 U36085 ( .A(n15967), .ZN(n11388) );
INV_X1 U36086 ( .A(n15966), .ZN(n11389) );
INV_X1 U36087 ( .A(n16124), .ZN(n11391) );
INV_X1 U36088 ( .A(n16118), .ZN(n11392) );
INV_X1 U36089 ( .A(n16046), .ZN(n11394) );
INV_X1 U36090 ( .A(n15972), .ZN(n11396) );
INV_X1 U36091 ( .A(n16045), .ZN(n11397) );
INV_X1 U36092 ( .A(n15971), .ZN(n11399) );
INV_X1 U36093 ( .A(n16116), .ZN(n11400) );
INV_X1 U36094 ( .A(n16117), .ZN(n11406) );
INV_X1 U36095 ( .A(n15812), .ZN(n11458) );
INV_X1 U36096 ( .A(n15803), .ZN(n11459) );
INV_X1 U36097 ( .A(n15793), .ZN(n11460) );
INV_X1 U36098 ( .A(crash_dump_o_96_), .ZN(n11464) );
INV_X1 U36099 ( .A(crash_dump_o_97_), .ZN(n11465) );
INV_X1 U36100 ( .A(crash_dump_o_101_), .ZN(n11466) );
INV_X1 U36101 ( .A(crash_dump_o_127_), .ZN(n11467) );
INV_X1 U36102 ( .A(n16132), .ZN(n11469) );
INV_X1 U36103 ( .A(n15929), .ZN(n11471) );
INV_X1 U36104 ( .A(n15927), .ZN(n11475) );
INV_X1 U36105 ( .A(cs_registers_i_mhpmcounter_0__3_), .ZN(n11478) );
INV_X1 U36106 ( .A(n15979), .ZN(n11509) );
INV_X1 U36107 ( .A(cs_registers_i_mhpmcounter_2__0_), .ZN(n11479) );
INV_X1 U36108 ( .A(n15926), .ZN(n11480) );
INV_X1 U36109 ( .A(n16047), .ZN(n11482) );
INV_X1 U36110 ( .A(n16129), .ZN(n11483) );
INV_X1 U36111 ( .A(crash_dump_o_65_), .ZN(n11485) );
INV_X1 U36112 ( .A(n16048), .ZN(n11488) );
INV_X1 U36113 ( .A(n16014), .ZN(n11489) );
INV_X1 U36114 ( .A(cs_registers_i_mhpmcounter_2__60_), .ZN(n11490) );
INV_X1 U36115 ( .A(cs_registers_i_mhpmcounter_2__29_), .ZN(n11491) );
INV_X1 U36116 ( .A(crash_dump_o_117_), .ZN(n11495) );
INV_X1 U36117 ( .A(crash_dump_o_85_), .ZN(n11496) );
INV_X1 U36118 ( .A(n16195), .ZN(n11499) );
INV_X1 U36119 ( .A(crash_dump_o_126_), .ZN(n11505) );
INV_X1 U36120 ( .A(crash_dump_o_94_), .ZN(n11506) );
INV_X1 U36121 ( .A(cs_registers_i_mhpmcounter_0__62_), .ZN(n11508) );
INV_X1 U36122 ( .A(cs_registers_i_mhpmcounter_0__31_), .ZN(n11510) );
INV_X1 U36123 ( .A(crash_dump_o_95_), .ZN(n11512) );
INV_X1 U36124 ( .A(crash_dump_o_69_), .ZN(n11513) );
endmodule